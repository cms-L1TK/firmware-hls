`timescale 1ns / 1ps

module SectorProcessor(
  input clk,
  input reset,
  input en_proc,
  input[2:0] bx_in_ProjectionRouter,
  output TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout,
  output TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout,
  output TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout,
  output TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout,
  output TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout,
  output TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout,
  output TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout,
  output TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb,
  output[7:0] TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr,
  input[59:0] TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout,
  input[7:0] TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout,
  input[7:0] TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout,
  output[2:0] bx_out_ProjectionRouter,
  output VMPROJ_L3PHIC20_dataarray_data_V_ena,
  output VMPROJ_L3PHIC20_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC20_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC20_dataarray_data_V_din,
  output VMPROJ_L3PHIC20_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC20_nentries_0_V_din,
  output VMPROJ_L3PHIC20_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC20_nentries_1_V_din,
  output VMPROJ_L3PHIC17_dataarray_data_V_ena,
  output VMPROJ_L3PHIC17_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC17_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC17_dataarray_data_V_din,
  output VMPROJ_L3PHIC17_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC17_nentries_0_V_din,
  output VMPROJ_L3PHIC17_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC17_nentries_1_V_din,
  output VMPROJ_L3PHIC22_dataarray_data_V_ena,
  output VMPROJ_L3PHIC22_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC22_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC22_dataarray_data_V_din,
  output VMPROJ_L3PHIC22_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC22_nentries_0_V_din,
  output VMPROJ_L3PHIC22_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC22_nentries_1_V_din,
  output VMPROJ_L3PHIC19_dataarray_data_V_ena,
  output VMPROJ_L3PHIC19_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC19_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC19_dataarray_data_V_din,
  output VMPROJ_L3PHIC19_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC19_nentries_0_V_din,
  output VMPROJ_L3PHIC19_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC19_nentries_1_V_din,
  output AP_L3PHIC_dataarray_data_V_ena,
  output AP_L3PHIC_dataarray_data_V_wea,
  output[9:0] AP_L3PHIC_dataarray_data_V_writeaddr,
  output[59:0] AP_L3PHIC_dataarray_data_V_din,
  output AP_L3PHIC_nentries_0_V_we,
  output[7:0] AP_L3PHIC_nentries_0_V_din,
  output AP_L3PHIC_nentries_1_V_we,
  output[7:0] AP_L3PHIC_nentries_1_V_din,
  output AP_L3PHIC_nentries_2_V_we,
  output[7:0] AP_L3PHIC_nentries_2_V_din,
  output AP_L3PHIC_nentries_3_V_we,
  output[7:0] AP_L3PHIC_nentries_3_V_din,
  output AP_L3PHIC_nentries_4_V_we,
  output[7:0] AP_L3PHIC_nentries_4_V_din,
  output AP_L3PHIC_nentries_5_V_we,
  output[7:0] AP_L3PHIC_nentries_5_V_din,
  output AP_L3PHIC_nentries_6_V_we,
  output[7:0] AP_L3PHIC_nentries_6_V_din,
  output AP_L3PHIC_nentries_7_V_we,
  output[7:0] AP_L3PHIC_nentries_7_V_din,
  output VMPROJ_L3PHIC24_dataarray_data_V_ena,
  output VMPROJ_L3PHIC24_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC24_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC24_dataarray_data_V_din,
  output VMPROJ_L3PHIC24_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC24_nentries_0_V_din,
  output VMPROJ_L3PHIC24_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC24_nentries_1_V_din,
  output VMPROJ_L3PHIC23_dataarray_data_V_ena,
  output VMPROJ_L3PHIC23_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC23_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC23_dataarray_data_V_din,
  output VMPROJ_L3PHIC23_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC23_nentries_0_V_din,
  output VMPROJ_L3PHIC23_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC23_nentries_1_V_din,
  output VMPROJ_L3PHIC18_dataarray_data_V_ena,
  output VMPROJ_L3PHIC18_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC18_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC18_dataarray_data_V_din,
  output VMPROJ_L3PHIC18_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC18_nentries_0_V_din,
  output VMPROJ_L3PHIC18_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC18_nentries_1_V_din,
  output VMPROJ_L3PHIC21_dataarray_data_V_ena,
  output VMPROJ_L3PHIC21_dataarray_data_V_wea,
  output[7:0] VMPROJ_L3PHIC21_dataarray_data_V_writeaddr,
  output[20:0] VMPROJ_L3PHIC21_dataarray_data_V_din,
  output VMPROJ_L3PHIC21_nentries_0_V_we,
  output[7:0] VMPROJ_L3PHIC21_nentries_0_V_din,
  output VMPROJ_L3PHIC21_nentries_1_V_we,
  output[7:0] VMPROJ_L3PHIC21_nentries_1_V_din,
  output ProjectionRouter_done
);

ProjectionRouter_BARRELPS_BARREL_8_3_0 PR_L3PHIC(
  .ap_clk(clk),
  .ap_rst(reset),
  .ap_start(en_proc),
  .ap_done(ProjectionRouter_done),
  .bx_V(bx_in_ProjectionRouter),
  .tproj1_dataarray_data_V_ce0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb),
  .tproj1_dataarray_data_V_address0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr),
  .tproj1_dataarray_data_V_q0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout),
  .tproj1_nentries_0_V(TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout),
  .tproj1_nentries_1_V(TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout),
  .tproj2_dataarray_data_V_ce0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb),
  .tproj2_dataarray_data_V_address0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr),
  .tproj2_dataarray_data_V_q0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout),
  .tproj2_nentries_0_V(TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout),
  .tproj2_nentries_1_V(TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout),
  .tproj3_dataarray_data_V_ce0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb),
  .tproj3_dataarray_data_V_address0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr),
  .tproj3_dataarray_data_V_q0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout),
  .tproj3_nentries_0_V(TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout),
  .tproj3_nentries_1_V(TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout),
  .tproj4_dataarray_data_V_ce0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb),
  .tproj4_dataarray_data_V_address0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr),
  .tproj4_dataarray_data_V_q0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout),
  .tproj4_nentries_0_V(TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout),
  .tproj4_nentries_1_V(TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout),
  .tproj5_dataarray_data_V_ce0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb),
  .tproj5_dataarray_data_V_address0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr),
  .tproj5_dataarray_data_V_q0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout),
  .tproj5_nentries_0_V(TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout),
  .tproj5_nentries_1_V(TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout),
  .tproj6_dataarray_data_V_ce0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb),
  .tproj6_dataarray_data_V_address0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr),
  .tproj6_dataarray_data_V_q0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout),
  .tproj6_nentries_0_V(TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout),
  .tproj6_nentries_1_V(TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout),
  .tproj7_dataarray_data_V_ce0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb),
  .tproj7_dataarray_data_V_address0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr),
  .tproj7_dataarray_data_V_q0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout),
  .tproj7_nentries_0_V(TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout),
  .tproj7_nentries_1_V(TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout),
  .tproj8_dataarray_data_V_ce0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb),
  .tproj8_dataarray_data_V_address0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr),
  .tproj8_dataarray_data_V_q0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout),
  .tproj8_nentries_0_V(TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout),
  .tproj8_nentries_1_V(TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout),
  .bx_o_V(bx_out_ProjectionRouter),
  .allproj_dataarray_data_V_ce0(AP_L3PHIC_dataarray_data_V_ena),
  .allproj_dataarray_data_V_we0(AP_L3PHIC_dataarray_data_V_wea),
  .allproj_dataarray_data_V_address0(AP_L3PHIC_dataarray_data_V_writeaddr),
  .allproj_dataarray_data_V_d0(AP_L3PHIC_dataarray_data_V_din),
  .allproj_nentries_0_V_ap_vld(AP_L3PHIC_nentries_0_V_we),
  .allproj_nentries_0_V(AP_L3PHIC_nentries_0_V_din),
  .allproj_nentries_1_V_ap_vld(AP_L3PHIC_nentries_1_V_we),
  .allproj_nentries_1_V(AP_L3PHIC_nentries_1_V_din),
  .allproj_nentries_2_V_ap_vld(AP_L3PHIC_nentries_2_V_we),
  .allproj_nentries_2_V(AP_L3PHIC_nentries_2_V_din),
  .allproj_nentries_3_V_ap_vld(AP_L3PHIC_nentries_3_V_we),
  .allproj_nentries_3_V(AP_L3PHIC_nentries_3_V_din),
  .allproj_nentries_4_V_ap_vld(AP_L3PHIC_nentries_4_V_we),
  .allproj_nentries_4_V(AP_L3PHIC_nentries_4_V_din),
  .allproj_nentries_5_V_ap_vld(AP_L3PHIC_nentries_5_V_we),
  .allproj_nentries_5_V(AP_L3PHIC_nentries_5_V_din),
  .allproj_nentries_6_V_ap_vld(AP_L3PHIC_nentries_6_V_we),
  .allproj_nentries_6_V(AP_L3PHIC_nentries_6_V_din),
  .allproj_nentries_7_V_ap_vld(AP_L3PHIC_nentries_7_V_we),
  .allproj_nentries_7_V(AP_L3PHIC_nentries_7_V_din),
  .vmproj1_dataarray_data_V_ce0(VMPROJ_L3PHIC17_dataarray_data_V_ena),
  .vmproj1_dataarray_data_V_we0(VMPROJ_L3PHIC17_dataarray_data_V_wea),
  .vmproj1_dataarray_data_V_address0(VMPROJ_L3PHIC17_dataarray_data_V_writeaddr),
  .vmproj1_dataarray_data_V_d0(VMPROJ_L3PHIC17_dataarray_data_V_din),
  .vmproj1_nentries_0_V_ap_vld(VMPROJ_L3PHIC17_nentries_0_V_we),
  .vmproj1_nentries_0_V(VMPROJ_L3PHIC17_nentries_0_V_din),
  .vmproj1_nentries_1_V_ap_vld(VMPROJ_L3PHIC17_nentries_1_V_we),
  .vmproj1_nentries_1_V(VMPROJ_L3PHIC17_nentries_1_V_din),
  .vmproj2_dataarray_data_V_ce0(VMPROJ_L3PHIC18_dataarray_data_V_ena),
  .vmproj2_dataarray_data_V_we0(VMPROJ_L3PHIC18_dataarray_data_V_wea),
  .vmproj2_dataarray_data_V_address0(VMPROJ_L3PHIC18_dataarray_data_V_writeaddr),
  .vmproj2_dataarray_data_V_d0(VMPROJ_L3PHIC18_dataarray_data_V_din),
  .vmproj2_nentries_0_V_ap_vld(VMPROJ_L3PHIC18_nentries_0_V_we),
  .vmproj2_nentries_0_V(VMPROJ_L3PHIC18_nentries_0_V_din),
  .vmproj2_nentries_1_V_ap_vld(VMPROJ_L3PHIC18_nentries_1_V_we),
  .vmproj2_nentries_1_V(VMPROJ_L3PHIC18_nentries_1_V_din),
  .vmproj3_dataarray_data_V_ce0(VMPROJ_L3PHIC19_dataarray_data_V_ena),
  .vmproj3_dataarray_data_V_we0(VMPROJ_L3PHIC19_dataarray_data_V_wea),
  .vmproj3_dataarray_data_V_address0(VMPROJ_L3PHIC19_dataarray_data_V_writeaddr),
  .vmproj3_dataarray_data_V_d0(VMPROJ_L3PHIC19_dataarray_data_V_din),
  .vmproj3_nentries_0_V_ap_vld(VMPROJ_L3PHIC19_nentries_0_V_we),
  .vmproj3_nentries_0_V(VMPROJ_L3PHIC19_nentries_0_V_din),
  .vmproj3_nentries_1_V_ap_vld(VMPROJ_L3PHIC19_nentries_1_V_we),
  .vmproj3_nentries_1_V(VMPROJ_L3PHIC19_nentries_1_V_din),
  .vmproj4_dataarray_data_V_ce0(VMPROJ_L3PHIC20_dataarray_data_V_ena),
  .vmproj4_dataarray_data_V_we0(VMPROJ_L3PHIC20_dataarray_data_V_wea),
  .vmproj4_dataarray_data_V_address0(VMPROJ_L3PHIC20_dataarray_data_V_writeaddr),
  .vmproj4_dataarray_data_V_d0(VMPROJ_L3PHIC20_dataarray_data_V_din),
  .vmproj4_nentries_0_V_ap_vld(VMPROJ_L3PHIC20_nentries_0_V_we),
  .vmproj4_nentries_0_V(VMPROJ_L3PHIC20_nentries_0_V_din),
  .vmproj4_nentries_1_V_ap_vld(VMPROJ_L3PHIC20_nentries_1_V_we),
  .vmproj4_nentries_1_V(VMPROJ_L3PHIC20_nentries_1_V_din),
  .vmproj5_dataarray_data_V_ce0(VMPROJ_L3PHIC21_dataarray_data_V_ena),
  .vmproj5_dataarray_data_V_we0(VMPROJ_L3PHIC21_dataarray_data_V_wea),
  .vmproj5_dataarray_data_V_address0(VMPROJ_L3PHIC21_dataarray_data_V_writeaddr),
  .vmproj5_dataarray_data_V_d0(VMPROJ_L3PHIC21_dataarray_data_V_din),
  .vmproj5_nentries_0_V_ap_vld(VMPROJ_L3PHIC21_nentries_0_V_we),
  .vmproj5_nentries_0_V(VMPROJ_L3PHIC21_nentries_0_V_din),
  .vmproj5_nentries_1_V_ap_vld(VMPROJ_L3PHIC21_nentries_1_V_we),
  .vmproj5_nentries_1_V(VMPROJ_L3PHIC21_nentries_1_V_din),
  .vmproj6_dataarray_data_V_ce0(VMPROJ_L3PHIC22_dataarray_data_V_ena),
  .vmproj6_dataarray_data_V_we0(VMPROJ_L3PHIC22_dataarray_data_V_wea),
  .vmproj6_dataarray_data_V_address0(VMPROJ_L3PHIC22_dataarray_data_V_writeaddr),
  .vmproj6_dataarray_data_V_d0(VMPROJ_L3PHIC22_dataarray_data_V_din),
  .vmproj6_nentries_0_V_ap_vld(VMPROJ_L3PHIC22_nentries_0_V_we),
  .vmproj6_nentries_0_V(VMPROJ_L3PHIC22_nentries_0_V_din),
  .vmproj6_nentries_1_V_ap_vld(VMPROJ_L3PHIC22_nentries_1_V_we),
  .vmproj6_nentries_1_V(VMPROJ_L3PHIC22_nentries_1_V_din),
  .vmproj7_dataarray_data_V_ce0(VMPROJ_L3PHIC23_dataarray_data_V_ena),
  .vmproj7_dataarray_data_V_we0(VMPROJ_L3PHIC23_dataarray_data_V_wea),
  .vmproj7_dataarray_data_V_address0(VMPROJ_L3PHIC23_dataarray_data_V_writeaddr),
  .vmproj7_dataarray_data_V_d0(VMPROJ_L3PHIC23_dataarray_data_V_din),
  .vmproj7_nentries_0_V_ap_vld(VMPROJ_L3PHIC23_nentries_0_V_we),
  .vmproj7_nentries_0_V(VMPROJ_L3PHIC23_nentries_0_V_din),
  .vmproj7_nentries_1_V_ap_vld(VMPROJ_L3PHIC23_nentries_1_V_we),
  .vmproj7_nentries_1_V(VMPROJ_L3PHIC23_nentries_1_V_din),
  .vmproj8_dataarray_data_V_ce0(VMPROJ_L3PHIC24_dataarray_data_V_ena),
  .vmproj8_dataarray_data_V_we0(VMPROJ_L3PHIC24_dataarray_data_V_wea),
  .vmproj8_dataarray_data_V_address0(VMPROJ_L3PHIC24_dataarray_data_V_writeaddr),
  .vmproj8_dataarray_data_V_d0(VMPROJ_L3PHIC24_dataarray_data_V_din),
  .vmproj8_nentries_0_V_ap_vld(VMPROJ_L3PHIC24_nentries_0_V_we),
  .vmproj8_nentries_0_V(VMPROJ_L3PHIC24_nentries_0_V_din),
  .vmproj8_nentries_1_V_ap_vld(VMPROJ_L3PHIC24_nentries_1_V_we),
  .vmproj8_nentries_1_V(VMPROJ_L3PHIC24_nentries_1_V_din)
);
endmodule
