--==========================================================================
-- CU Boulder
-------------------------------------------------------------------------------
--! @file
--! @brief Test bench for the track finding top using TextIO.
--! @author Robert Glein
--! @date 2020-05-18
--! @version v.1.0
--=============================================================================

--! Standard library
library ieee;
--! Standard package
use ieee.std_logic_1164.all;
--! Signed/unsigned calculations
use ieee.numeric_std.all;
--! Math real
use ieee.math_real.all;
--! TextIO
use ieee.std_logic_textio.all;
--! Standard functions
library std;
--! Standard TextIO functions
use std.textio.all;

--! Xilinx library
library unisim;
--! Xilinx package
use unisim.vcomponents.all;

--! User packages
use work.mytypes_pkg.all;



--! @brief TB
entity tb_top_tf is
end tb_top_tf;

--! @brief TB
architecture behavior of tb_top_tf is
  -- ########################### Types ###########################
  type t_str_array_TPROJ is array(natural range <>) of string(1 to 103); --! String array
  type t_str_array_VMSME is array(natural range <>) of string(1 to 79);  --! String array
  type t_str_array_VMP   is array(natural range <>) of string(1 to 41);  --! String array
  type t_str_array_CM    is array(natural range <>) of string(1 to 37);  --! String array
  type t_str_array_FM    is array(natural range <>) of string(1 to 42);  --! String array
  type t_myarray_1d_1d_int    is array(natural range <>) of t_myarray_1d_int(0 to MAX_EVENTS-1);                      --! 1x1D array of int
  type t_myarray_1d_2d_int    is array(natural range <>) of t_myarray_2d_int(0 to MAX_EVENTS-1,0 to N_MEM_BINS-1);    --! 1x2D array of int
  type t_myarray_1d_2d_slv_2p is array(natural range <>) of t_myarray_2d_slv(0 to MAX_EVENTS-1,0 to 2*PAGE_OFFSET-1); --! 1x2D array of slv
  type t_myarray_1d_2d_slv_8p is array(natural range <>) of t_myarray_2d_slv(0 to MAX_EVENTS-1,0 to 8*PAGE_OFFSET-1); --! 1x2D array of slv

  -- ########################### Constant Definitions ###########################
  -- ############ Please change the constants in this section ###################
  constant N_ME_IN_CHAIN     : integer := 8; --! Number of match engines in chain
  constant INST_TOP_TF       : integer := 2;          --! Instantiate top_tf or others
                                                      --! 0: Generated prmemc chain
                                                      --! 1: top_tf
                                                      --! 2: top_tf_full
  constant CLK_PERIOD        : time    := 4.16667 ns; --! 240 MHz
  constant DEBUG             : boolean := true;       --! Debug off/on
  constant VMSME_DELAY       : integer := 1-1;        --! Number of BX delays (can be written early 8 pages)
  constant AS_DELAY          : integer := 2-1;        --! Number of BX delays (can be written early 8 pages)
  constant MEM_READ_DELAY    : integer := 2;          --! Number of memory read delay
  constant FILE_IN_TPROJ : t_str_array_TPROJ(0 to N_ME_IN_CHAIN-1) := ("../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L1L2F_L3PHIC_04.dat", --! Input files
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L1L2G_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L1L2H_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L1L2I_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L1L2J_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L5L6B_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L5L6C_L3PHIC_04.dat",
                                                                       "../../../../../../../emData/MemPrints/TrackletProjections/TrackletProjections_TPROJ_L5L6D_L3PHIC_04.dat" );
  constant FILE_IN_VMSME : t_str_array_VMSME(0 to N_ME_IN_CHAIN-1) := ("../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC17n1_04.dat", --! Input files
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC18n1_04.dat",
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC19n1_04.dat",
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC20n1_04.dat", -- Used by lastest ME HLS c(o)sim
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC21n1_04.dat",
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC22n1_04.dat",
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC23n1_04.dat",
                                                                       "../../../../../../../emData/MemPrints/VMStubsME/VMStubs_VMSME_L3PHIC24n1_04.dat" );
  constant FILE_IN_AS        : string := "../../../../../../../emData/MemPrints/Stubs/AllStubs_AS_L3PHICn6_04.dat"; --! Input file
  constant FILE_OUT_VMP      : t_str_array_VMP(0 to N_ME_IN_CHAIN-1) := ("../../../../../TextIO/VMPROJ_L3PHIC17.txt", --! Output file for VMP
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC18.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC19.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC20.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC21.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC22.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC23.txt",
                                                                         "../../../../../TextIO/VMPROJ_L3PHIC24.txt" );
  constant FILE_OUT_AP       : string := "../../../../../TextIO/AP_L3PHIC.txt";  --! Output file for AP
  constant FILE_OUT_CM       : t_str_array_CM(0 to N_ME_IN_CHAIN-1) :=  ("../../../../../TextIO/CM_L3PHIC17.txt", --! Output file for CM
                                                                         "../../../../../TextIO/CM_L3PHIC18.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC19.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC20.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC21.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC22.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC23.txt",
                                                                         "../../../../../TextIO/CM_L3PHIC24.txt" );
  constant FILE_OUT_FM       : t_str_array_FM(0 to 1) :=  ("../../../../../TextIO/FM_L1L2XX_L3PHIC.txt", --! Output file for FM
                                                           "../../../../../TextIO/FM_L5L6XX_L3PHIC.txt" );

  -- ########################### Signals ###########################
  -- ### UUT signals ###
  signal clk       : std_logic := '0';
  signal reset     : std_logic := '1';
  signal PR_start  : std_logic := '0';
  signal PR_idle   : std_logic;
  signal PR_ready  : std_logic;
  signal PR_bx_in  : std_logic_vector(2 downto 0) := (others => '0');
  -- For TrackletProjections memories
  signal TPROJ_L3PHIC_dataarray_data_V_wea       : t_myarray8_1b   := (others => '0');
  signal TPROJ_L3PHIC_dataarray_data_V_writeaddr : t_myarray8_8b   := (others => (others => '0'));
  signal TPROJ_L3PHIC_dataarray_data_V_din       : t_myarray8_60b  := (others => (others => '0'));
  signal TPROJ_L3PHIC_nentries_V_we  : t_myarray2_8_1b := (others => (others => '0'));
  signal TPROJ_L3PHIC_nentries_V_din : t_myarray2_8_8b := (others => (others => (others => '0')));
  -- For VMStubME memories
  signal VMSME_L3PHIC17to24n1_dataarray_data_V_wea       : t_myarray8_1b  := (others => '0');
  signal VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr : t_myarray8_10b  := (others => (others => '0'));
  signal VMSME_L3PHIC17to24n1_dataarray_data_V_din       : t_myarray8_14b := (others => (others => '0'));
  signal VMSME_L3PHIC17to24n1_nentries_V_we  : t_myarray8_8_8_1b := (others => (others => (others => '0')));             -- (#page, #bin, #mem)
  signal VMSME_L3PHIC17to24n1_nentries_V_din : t_myarray8_8_8_4b := (others => (others => (others => (others => '0')))); -- (#page, #bin, #mem)
  -- For AllStubs memories
  signal AS_L3PHICn4_dataarray_data_V_wea       : std_logic                     := '0';
  signal AS_L3PHICn4_dataarray_data_V_writeaddr : std_logic_vector(9 downto 0)  := (others => '0');
  signal AS_L3PHICn4_dataarray_data_V_din       : std_logic_vector(35 downto 0) := (others => '0');
  signal AS_L3PHICn4_nentries_V_we  : t_myarray8_1b := (others => '0');
  signal AS_L3PHICn4_nentries_V_din : t_myarray8_8b := (others => (others => '0'));
  -- FullMatches output
  signal FM_L1L2XX_L3PHIC_dataarray_data_V_enb      : std_logic                     := '0';
  signal FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0)  := (others => '0');
  signal FM_L1L2XX_L3PHIC_dataarray_data_V_dout     : std_logic_vector(44 downto 0);
  signal FM_L1L2XX_L3PHIC_nentries_V_dout : t_myarray2_8b;
  signal FM_L5L6XX_L3PHIC_dataarray_data_V_enb      : std_logic                     := '0';
  signal FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0)  := (others => '0');
  signal FM_L5L6XX_L3PHIC_dataarray_data_V_dout     : std_logic_vector(44 downto 0);
  signal FM_L5L6XX_L3PHIC_nentries_V_dout : t_myarray2_8b;
  -- MatchCalculator outputs
  signal MC_bx_out     : std_logic_vector(2 downto 0);
  signal MC_bx_out_vld : std_logic;
  signal MC_done       : std_logic;
  -- ### Other signals ###
  signal PR_start_tmp                       : std_logic := '0';
  signal TPROJ_L3PHICn4_data_arr            : t_myarray_1d_2d_slv_2p(0 to N_ME_IN_CHAIN-1);
  signal TPROJ_L3PHICn4_n_entries_arr       : t_myarray_1d_1d_int(0 to N_ME_IN_CHAIN-1);
  signal VMSME_L3PHIC17to24n1_data_arr      : t_myarray_1d_2d_slv_8p(0 to N_ME_IN_CHAIN-1);
  signal VMSME_L3PHIC17to24n1_n_entries_arr : t_myarray_1d_2d_int(0 to N_ME_IN_CHAIN-1);
  signal AS_L3PHICn4_data_arr               : t_myarray_2d_slv(0 to MAX_EVENTS-1,0 to 8*PAGE_OFFSET-1);
  signal AS_L3PHICn4_n_entries_arr          : t_myarray_1d_int(0 to MAX_EVENTS-1);
  signal bx_cnt                             : integer := 0; -- BX counter
  signal page_cnt2                          : integer := 0; -- Page counter
  signal page_cnt8                          : integer := 0; -- Page counter
  -- ### Signals for top_tf_full only (VHDL does not support conditional signal declaration) ###
  -- ProjectionRouter outputs
  signal PR_done       : std_logic := '0';
  signal PR_bx_out     : std_logic_vector(2 downto 0);
  signal PR_bx_out_vld : std_logic;
  -- AllProjection output
  signal AP_L3PHIC_dataarray_data_V_wea       : std_logic;
  signal AP_L3PHIC_dataarray_data_V_writeaddr : std_logic_vector(9 downto 0);
  signal AP_L3PHIC_dataarray_data_V_din       : std_logic_vector(59 downto 0);
  --signal AP_L3PHIC_nentries_V_we  : t_myarray8_1b;
  --signal AP_L3PHIC_nentries_V_din : t_myarray8_8b;
  -- VMProjection output
  signal VMPROJ_L3PHIC17to24_dataarray_data_V_wea       : t_myarray8_1b;
  signal VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr : t_myarray8_8b;
  signal VMPROJ_L3PHIC17to24_dataarray_data_V_din       : t_myarray8_21b;
  --signal VMPROJ_L3PHIC17to24_nentries_V_we  : t_myarray2_8_1b;
  --signal VMPROJ_L3PHIC17to24_nentries_V_din : t_myarray2_8_8b;
  -- MatchEngine output
  signal ME_bx_out     : t_myarray8_3b;
  signal ME_bx_out_vld : t_myarray8_1b;
  signal ME_all_done   : std_logic := '0';
  -- CandidateMatch output
  signal CM_L3PHIC17to24_dataarray_data_V_wea       : t_myarray8_1b;
  signal CM_L3PHIC17to24_dataarray_data_V_writeaddr : t_myarray8_8b;
  signal CM_L3PHIC17to24_dataarray_data_V_din       : t_myarray8_14b;
  --signal CM_L3PHIC17to24_nentries_V_we  : t_myarray2_8_1b;
  --signal CM_L3PHIC17to24_nentries_V_din : t_myarray2_8_8b;


begin

  -- ########################### Processes ###########################

  --! @brief Clock process ---------------------------------------
  CLK_process : process
  begin
    clk <= '1';
    wait for CLK_PERIOD/2;
    clk <= '0';
    wait for CLK_PERIOD/2;
  end process CLK_process;

  --! @brief Read emData process ---------------------------------------
  read_data : process
    variable v_TPROJ_L3PHICn4_data_arr            : t_myarray_1d_2d_slv_2p(0 to N_ME_IN_CHAIN-1);
    variable v_TPROJ_L3PHICn4_n_entries_arr       : t_myarray_1d_1d_int(0 to N_ME_IN_CHAIN-1);
    variable v_VMSME_L3PHIC17to24n1_data_arr      : t_myarray_1d_2d_slv_8p(0 to N_ME_IN_CHAIN-1);
    variable v_VMSME_L3PHIC17to24n1_n_entries_arr : t_myarray_1d_2d_int(0 to N_ME_IN_CHAIN-1);
    variable v_AS_L3PHICn4_data_arr               : t_myarray_2d_slv(0 to MAX_EVENTS-1,0 to N_ME_IN_CHAIN*PAGE_OFFSET-1);
    variable v_AS_L3PHICn4_n_entries_arr          : t_myarray_1d_int(0 to MAX_EVENTS-1);
    variable v_line_in : line; -- Line for debug
  begin
    -- TPROJ
    l_TPROJ_read : for i in 0 to N_ME_IN_CHAIN-1 loop
      read_emData_2p (FILE_IN_TPROJ(i), v_TPROJ_L3PHICn4_data_arr(i), v_TPROJ_L3PHICn4_n_entries_arr(i));
      if DEBUG=true then write(v_line_in, string'("TPROJ_i: ")); write(v_line_in, i); write(v_line_in, string'(";   v_TPROJ_L3PHICn4_data_arr(i)(0,0): ")); hwrite(v_line_in, v_TPROJ_L3PHICn4_data_arr(i)(0,0)); writeline(output, v_line_in); end if;
      if DEBUG=true then write(v_line_in, string'("TPROJ_i: ")); write(v_line_in, i); write(v_line_in, string'(";   v_TPROJ_L3PHICn4_n_entries_arr(i)(0): ")); write(v_line_in, v_TPROJ_L3PHICn4_n_entries_arr(i)(0)); writeline(output, v_line_in); end if;
    end loop l_TPROJ_read;
    if DEBUG=true then write(v_line_in, string'("v_TPROJ_L3PHICn4_data_arr(0)(99,0+128): ")); hwrite(v_line_in, v_TPROJ_L3PHICn4_data_arr(0)(99,0+128)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_TPROJ_L3PHICn4_data_arr(0)(99,3+128): ")); hwrite(v_line_in, v_TPROJ_L3PHICn4_data_arr(0)(99,3+128)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_TPROJ_L3PHICn4_n_entries_arr(0)(99): "));   write(v_line_in, v_TPROJ_L3PHICn4_n_entries_arr(0)(99)); writeline(output, v_line_in); end if;
    -- VMSME
    l_VMSME_read : for i in 0 to N_ME_IN_CHAIN-1 loop
      read_emData_8p_bin (FILE_IN_VMSME(i), v_VMSME_L3PHIC17to24n1_data_arr(i), v_VMSME_L3PHIC17to24n1_n_entries_arr(i));
      if DEBUG=true then write(v_line_in, string'("VMSME_i: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_data_arr(i)(0,0): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(i)(0,0)); writeline(output, v_line_in); end if;
      if DEBUG=true then write(v_line_in, string'("VMSME_i: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_n_entries_arr(i)(0,0): ")); write(v_line_in, v_VMSME_L3PHIC17to24n1_n_entries_arr(i)(0,0)); writeline(output, v_line_in); end if;
    end loop l_VMSME_read;
    if DEBUG=true then write(v_line_in, string'("v_VMSME_L3PHIC17to24n1_data_arr(0)(99,3*PAGE_OFFSET+7*N_ENTRIES_PER_MEM_BINS): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(0)(99,3*PAGE_OFFSET+7*N_ENTRIES_PER_MEM_BINS)); writeline(output, v_line_in); end if;
      if DEBUG=true then write(v_line_in, string'("v_VMSME_L3PHIC17to24n1_n_entries_arr(0)(99,7): ")); write(v_line_in, v_VMSME_L3PHIC17to24n1_n_entries_arr(0)(99,7)); writeline(output, v_line_in); end if;
    l_VMSME_debug0 : for i in 0 to 64 loop -- until last utilized addr
      if DEBUG=true then write(v_line_in, string'("addr: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_data_arr(0)(0,addr): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(0)(0,i)); writeline(output, v_line_in); end if;
    end loop l_VMSME_debug0;
    l_VMSME_debug9 : for i in 1*PAGE_OFFSET to 1*PAGE_OFFSET+(5*16+1) loop -- until last utilized addr
      if DEBUG=true then write(v_line_in, string'("addr: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_data_arr(6)(9,addr): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(6)(9,i)); writeline(output, v_line_in); end if;
    end loop l_VMSME_debug9;
    l_VMSME_debug23 : for i in 7*PAGE_OFFSET to 7*PAGE_OFFSET+(6*16+4) loop -- until last utilized addr
      if DEBUG=true then write(v_line_in, string'("addr: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_data_arr(4)(23,addr): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(4)(23,i)); writeline(output, v_line_in); end if;
    end loop l_VMSME_debug23;
    l_VMSME_debug99 : for i in 3*PAGE_OFFSET to 3*PAGE_OFFSET+(7*16) loop -- until last utilized addr
      if DEBUG=true then write(v_line_in, string'("addr: ")); write(v_line_in, i); write(v_line_in, string'(";   v_VMSME_L3PHIC17to24n1_data_arr(0)(99,addr): ")); hwrite(v_line_in, v_VMSME_L3PHIC17to24n1_data_arr(0)(99,i)); writeline(output, v_line_in); end if;
    end loop l_VMSME_debug99;
    -- AS
    read_emData_8p (FILE_IN_AS, v_AS_L3PHICn4_data_arr, v_AS_L3PHICn4_n_entries_arr);
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_data_arr(0,0): "));         hwrite(v_line_in, v_AS_L3PHICn4_data_arr(0,0)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_data_arr(0,71): "));        hwrite(v_line_in, v_AS_L3PHICn4_data_arr(0,71)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_n_entries_arr(0): "));       write(v_line_in, v_AS_L3PHICn4_n_entries_arr(0)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_data_arr(99,0+128*3): "));  hwrite(v_line_in, v_AS_L3PHICn4_data_arr(99,0+128*3)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_data_arr(99,35+128*3): ")); hwrite(v_line_in, v_AS_L3PHICn4_data_arr(99,35+128*3)); writeline(output, v_line_in); end if;
    if DEBUG=true then write(v_line_in, string'("v_AS_L3PHICn4_n_entries_arr(99): "));      write(v_line_in, v_AS_L3PHICn4_n_entries_arr(99)); writeline(output, v_line_in); end if;
    -- Map variables to signals
    TPROJ_L3PHICn4_data_arr            <= v_TPROJ_L3PHICn4_data_arr;
    TPROJ_L3PHICn4_n_entries_arr       <= v_TPROJ_L3PHICn4_n_entries_arr;
    VMSME_L3PHIC17to24n1_data_arr      <= v_VMSME_L3PHIC17to24n1_data_arr;
    VMSME_L3PHIC17to24n1_n_entries_arr <= v_VMSME_L3PHIC17to24n1_n_entries_arr;
    AS_L3PHICn4_data_arr               <= v_AS_L3PHICn4_data_arr;
    AS_L3PHICn4_n_entries_arr          <= v_AS_L3PHICn4_n_entries_arr;
    wait;
  end process read_data;

  --! @brief Playback process ---------------------------------------
  --! @BoBX0: en_proc=0,   w TPROJ p1,
  --! @BoBX1: en_proc=1,   w TPROJ p2,  w VMSME p1
  --! @BoBX2: en_proc=1,   w TPROJ p1,  w VMSME p2, w AS p1
  --! @BoBX3: en_proc=1,   w TPROJ p2,  w VMSME p3, w AS p2
  --! @BoBX3: en_proc=1,   w TPROJ p1,  w VMSME p4, w AS p3
  --! ...
  playback : process
    variable v_page_cnt2_d0            : integer := 0; -- Page counter 
    variable v_page_cnt2_d1            : integer := 0; -- Page counter delayed by one
    variable v_page_cnt8               : integer := 0; -- Page counter
    variable v_VMSME_n_entries_bin     : t_myarray_1d_int(0 to N_ME_IN_CHAIN-1) := (others => 0); -- Number of VMSME entries per bin
    variable v_VMSME_n_entries_bin_cnt : t_myarray_1d_int(0 to N_ME_IN_CHAIN-1) := (others => 0); -- Counter of VMSME entries per bin
    variable v_bin_cnt                 : t_myarray_1d_int(0 to N_ME_IN_CHAIN-1) := (others => 0); -- Bin counter
    variable v_last_bin                : boolean := false; -- Last bin tag
    variable v_line_in : line; -- Line for debug
  begin
    wait for CLK_PERIOD; -- Let the read process finish
    reset <= '0';           -- Reset cycle
    l_BX : for v_bx_cnt in -1 to MAX_EVENTS+10 loop -- -1 (to write the first memories before starting) to 110 (+10 to let later modules and write finish)
      bx_cnt         <= v_bx_cnt;       -- Update the signal
      v_page_cnt2_d0 := v_bx_cnt mod 2;          -- mod 2
      v_page_cnt2_d1 := (v_bx_cnt+1) mod 2;      -- mod 2
      v_page_cnt8    := v_bx_cnt mod N_MEM_BINS; -- mod 8
      page_cnt2      <= v_page_cnt2_d0; -- Update the signal
      page_cnt8      <= v_page_cnt8;    -- Update the signal
      v_bin_cnt      := (others => 0);
      v_VMSME_n_entries_bin_cnt := (others => 0);
      PR_bx_in <= std_logic_vector(to_unsigned(v_bx_cnt, PR_bx_in'length));
      l_addr : for addr in 0 to MAX_ENTRIES-1 loop -- 0 to 107
        l_copies : for cp in 0 to N_ME_IN_CHAIN-1 loop -- 0 to 7 -- Unable to assign arrays directly
          v_last_bin := false; -- Default assigment
          -- TPROJ
          if (v_bx_cnt<MAX_EVENTS-1) then -- Start early
            TPROJ_L3PHIC_dataarray_data_V_wea <= (others => '1');
            TPROJ_L3PHIC_nentries_V_we        <= (others => (others => '1'));
            TPROJ_L3PHIC_dataarray_data_V_writeaddr(cp) <= std_logic_vector(to_unsigned(addr+PAGE_OFFSET*v_page_cnt2_d1, TPROJ_L3PHIC_dataarray_data_V_writeaddr(0)'length));
            TPROJ_L3PHIC_dataarray_data_V_din(cp)       <= TPROJ_L3PHICn4_data_arr(cp)(v_bx_cnt+1,addr+PAGE_OFFSET*v_page_cnt2_d1) (TPROJ_L3PHIC_dataarray_data_V_din(0)'length-1 downto 0);
            TPROJ_L3PHIC_nentries_V_din(v_page_cnt2_d1)(cp) <= std_logic_vector(to_unsigned(TPROJ_L3PHICn4_n_entries_arr(cp)(v_bx_cnt+1), TPROJ_L3PHIC_nentries_V_din(0)(0)'length));
          end if;
          -- VMSME & PR_start
          PR_start <= '0'; -- Default assigment
          if (v_bx_cnt>=VMSME_DELAY and v_bx_cnt<MAX_EVENTS-1) then -- Start after delay of BXs
            if (PR_ready='1' or PR_idle='1') and PR_start_tmp='0' then -- Control PR start
              PR_start_tmp <= '1';
            else
              PR_start_tmp <= '0';
            end if;
            PR_start <= PR_start_tmp;
            VMSME_L3PHIC17to24n1_dataarray_data_V_wea(cp) <= '1';                                     -- Default assigment
            VMSME_L3PHIC17to24n1_nentries_V_we            <= (others => (others => (others => '1'))); -- Default assigment
            if v_bin_cnt(cp)<=N_MEM_BINS-1 then -- Valid bin
              v_VMSME_n_entries_bin(cp) := VMSME_L3PHIC17to24n1_n_entries_arr(cp)(v_bx_cnt-VMSME_DELAY,v_bin_cnt(cp));
              VMSME_L3PHIC17to24n1_nentries_V_din(((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS))(v_bin_cnt(cp))(cp) <= std_logic_vector(to_unsigned(v_VMSME_n_entries_bin(cp), VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(0)'length));
            end if;
            l_bin_empty : while (v_VMSME_n_entries_bin(cp)<=0) loop -- Bin empty
              v_bin_cnt(cp)             := v_bin_cnt(cp) +1; -- Skip empty bin
              if v_bin_cnt(cp)<=N_MEM_BINS-1 then -- Valid bin
                v_VMSME_n_entries_bin(cp) := VMSME_L3PHIC17to24n1_n_entries_arr(cp)(v_bx_cnt-VMSME_DELAY,v_bin_cnt(cp));
                VMSME_L3PHIC17to24n1_nentries_V_din(((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS))(v_bin_cnt(cp))(cp) <= std_logic_vector(to_unsigned(v_VMSME_n_entries_bin(cp), VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(0)'length));
              else
                v_bin_cnt(cp) := N_MEM_BINS;
                exit;
              end if;
            end loop l_bin_empty;
            if v_bin_cnt(cp)<=N_MEM_BINS-1 then -- Valid bin
              VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(cp) <=                            std_logic_vector(to_unsigned((v_bin_cnt(cp)*N_ENTRIES_PER_MEM_BINS+v_VMSME_n_entries_bin_cnt(cp)) + (PAGE_OFFSET*((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS)), VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(0)'length));
              VMSME_L3PHIC17to24n1_dataarray_data_V_din(cp)       <= VMSME_L3PHIC17to24n1_data_arr(cp)(v_bx_cnt-VMSME_DELAY, (v_bin_cnt(cp)*N_ENTRIES_PER_MEM_BINS+v_VMSME_n_entries_bin_cnt(cp)) + (PAGE_OFFSET*((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS))) (VMSME_L3PHIC17to24n1_dataarray_data_V_din(0)'length-1 downto 0);
              if (DEBUG=true and ((v_bx_cnt=9 and cp=6) or (v_bx_cnt=23 and cp=4))) then write(v_line_in, string'("v_bx_cnt: ")); write(v_line_in, v_bx_cnt); write(v_line_in, string'(";   cp: ")); write(v_line_in, cp); writeline(output, v_line_in); end if;
              if (DEBUG=true and ((v_bx_cnt=9 and cp=6) or (v_bx_cnt=23 and cp=4))) then write(v_line_in, string'("VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(cp): ")); write(v_line_in, ((v_bin_cnt(cp)*N_ENTRIES_PER_MEM_BINS+v_VMSME_n_entries_bin_cnt(cp)) + (PAGE_OFFSET*((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS)))); writeline(output, v_line_in); end if;
              if (DEBUG=true and ((v_bx_cnt=9 and cp=6) or (v_bx_cnt=23 and cp=4))) then write(v_line_in, string'("VMSME_L3PHIC17to24n1_dataarray_data_V_din(cp): ")); hwrite(v_line_in, VMSME_L3PHIC17to24n1_data_arr(cp)(v_bx_cnt-VMSME_DELAY, (v_bin_cnt(cp)*N_ENTRIES_PER_MEM_BINS+v_VMSME_n_entries_bin_cnt(cp)) + (PAGE_OFFSET*((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS))) (VMSME_L3PHIC17to24n1_dataarray_data_V_din(0)'length-1 downto 0)); writeline(output, v_line_in); end if;
              if (DEBUG=true and ((v_bx_cnt=9 and cp=6) or (v_bx_cnt=23 and cp=4))) then write(v_line_in, string'("v_VMSME_n_entries_bin_cnt(cp): ")); write(v_line_in, v_VMSME_n_entries_bin_cnt(cp)); write(v_line_in, string'(";   v_VMSME_n_entries_bin(cp): ")); write(v_line_in, v_VMSME_n_entries_bin(cp)); write(v_line_in, string'(";   v_bin_cnt(cp): ")); write(v_line_in, v_bin_cnt(cp)); writeline(output, v_line_in); end if;
            end if;
            --if DEBUG=true then assert (addr>1 or v_bx_cnt>0) report "addr = " & integer'image(addr) & ";   cp = " & integer'image(addr) & ";   v_bin_cnt(0) = " & integer'image(v_bin_cnt(0)) & ";   v_VMSME_n_entries_bin_cnt(cp) = " & integer'image(v_VMSME_n_entries_bin_cnt(cp)) & ";   waddr = " & integer'image((v_bin_cnt(0)*N_ENTRIES_PER_MEM_BINS+v_VMSME_n_entries_bin_cnt(cp)) + (PAGE_OFFSET*((v_page_cnt8-VMSME_DELAY) mod N_MEM_BINS))) severity note; end if;
            if v_VMSME_n_entries_bin_cnt(cp)>=v_VMSME_n_entries_bin(cp)-1 then -- End of bin entries
              if (v_bin_cnt(cp)=N_MEM_BINS-1) then -- Last bin
                v_last_bin := true;
              end if;
              v_bin_cnt(cp)                 := v_bin_cnt(cp) +1;
              v_VMSME_n_entries_bin_cnt(cp) := 0;
              if (v_bin_cnt(cp)>=N_MEM_BINS) then
                v_bin_cnt(cp)               := N_MEM_BINS; -- End of write for this addr
              end if;
            else
              v_VMSME_n_entries_bin_cnt(cp) := v_VMSME_n_entries_bin_cnt(cp) +1;
            end if;
            if v_bin_cnt(cp)>N_MEM_BINS-1 then -- Invalid bin
              v_bin_cnt(cp) := N_MEM_BINS; 
              if v_last_bin=false then
                VMSME_L3PHIC17to24n1_dataarray_data_V_wea(cp) <= '0';
                VMSME_L3PHIC17to24n1_nentries_V_we            <= (others => (others => (others => '0')));
              end if;
            end if;
          end if;
          -- AS
          if (v_bx_cnt>=AS_DELAY and v_bx_cnt<MAX_EVENTS-1) then -- Start after delay of BXs
            AS_L3PHICn4_dataarray_data_V_wea <= '1';
            AS_L3PHICn4_nentries_V_we        <= (others => '1');
            AS_L3PHICn4_dataarray_data_V_writeaddr  <= std_logic_vector(to_unsigned(addr+(PAGE_OFFSET*((v_page_cnt8-AS_DELAY) mod N_MEM_BINS)),AS_L3PHICn4_dataarray_data_V_writeaddr'length));
            AS_L3PHICn4_dataarray_data_V_din        <= AS_L3PHICn4_data_arr(v_bx_cnt-AS_DELAY,addr+(PAGE_OFFSET*((v_page_cnt8-AS_DELAY) mod N_MEM_BINS))) (AS_L3PHICn4_dataarray_data_V_din'length-1 downto 0); 
            AS_L3PHICn4_nentries_V_din((v_page_cnt8-AS_DELAY) mod N_MEM_BINS) <= std_logic_vector(to_unsigned(AS_L3PHICn4_n_entries_arr(v_bx_cnt-AS_DELAY), AS_L3PHICn4_nentries_V_din(0)'length));
          end if;
        end loop l_copies;
        wait for CLK_PERIOD; -- Main time control
        --if DEBUG=true then assert (v_bx_cnt>0) report "addr = " & integer'image(addr) & ";   VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(0) = " & integer'image(to_integer(unsigned(VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(0)))) severity note; end if;
      end loop l_addr;
    end loop l_BX;
    wait for CLK_PERIOD;
  end process playback;

  --! @brief TextIO process for writting the output ---------------------------------------
  write_result : process
    file     file_out_L1L2 : text open WRITE_MODE is FILE_OUT_FM(0); -- Text - a file of character strings
    file     file_out_L5L6 : text open WRITE_MODE is FILE_OUT_FM(1); -- Text - a file of character strings
    variable v_line   : line;                                        -- Line - one string from a text
    variable v_FM_L1L2XX_L3PHIC_dataarray_data_V_enb_d : std_logic_vector(MEM_READ_DELAY-1 downto 0) := (others => '0'); -- Delay vector
    variable v_FM_L5L6XX_L3PHIC_dataarray_data_V_enb_d : std_logic_vector(MEM_READ_DELAY-1 downto 0) := (others => '0'); -- Delay vector
  begin
    -- Write file header
    write(v_line, string'("time"), right, 20); write(v_line, string'("BX#"), right, 4);
    write(v_line, string'("reset"), right, 6);
    write(v_line, string'("n_ent_p0"), right, 9); write(v_line, string'("n_ent_p1"), right, 9); write(v_line, string'("enb"), right, 4);
    write(v_line, string'("readaddr"), right, 9);  write(v_line, string'("FM_L1L2XX_L3PHIC_dataarray_data_V_dout"), right, 39);
    write(v_line, string'("MC_done"), right, 9);  write(v_line, string'("MC_bx_out_vld"), right, 14); write(v_line, string'("MC_bx_out"), right, 10);
    writeline (file_out_L1L2, v_line); -- Write line
    write(v_line, string'("time"), right, 20); write(v_line, string'("BX#"), right, 4);
    write(v_line, string'("reset"), right, 6);
    write(v_line, string'("n_ent_p0"), right, 9); write(v_line, string'("n_ent_p1"), right, 9); write(v_line, string'("enb"), right, 4);
    write(v_line, string'("readaddr"), right, 9);  write(v_line, string'("FM_L5L6XX_L3PHIC_dataarray_data_V_dout"), right, 39);
    write(v_line, string'("MC_done"), right, 9);  write(v_line, string'("MC_bx_out_vld"), right, 14); write(v_line, string'("MC_bx_out"), right, 10);
    writeline (file_out_L5L6, v_line); -- Write line
    wait until rising_edge(MC_done); -- Wait for first result
    l_BX : for v_bx_cnt in 0 to MAX_EVENTS-1 loop -- 0 to 99
      l_addr : for addr in 0 to MAX_ENTRIES-1+MEM_READ_DELAY loop -- 0 to 109
        if (addr <= MAX_ENTRIES-1) then -- w/o MEM_READ_DELAY
-- todo: write all 256 addr to file; pause playback and en_proc (wait for readout done)
          if (v_bx_cnt mod 2)=0 then -- 1. page
            if (addr < (to_integer(unsigned(FM_L1L2XX_L3PHIC_nentries_V_dout(0))))) then -- Only read number of entries: Switch off in complete read out mode
              FM_L1L2XX_L3PHIC_dataarray_data_V_enb <= '1';
            else
              FM_L1L2XX_L3PHIC_dataarray_data_V_enb <= '0';
            end if;
            if (addr < (to_integer(unsigned(FM_L5L6XX_L3PHIC_nentries_V_dout(0))))) then -- Only read number of entries: Switch off in complete read out mode
              FM_L5L6XX_L3PHIC_dataarray_data_V_enb <= '1';
            else
              FM_L5L6XX_L3PHIC_dataarray_data_V_enb <= '0';
            end if;
          else                       -- 2. page
            if (addr < (to_integer(unsigned(FM_L1L2XX_L3PHIC_nentries_V_dout(1))))) then -- Only read number of entries: Switch off in complete read out mode
              FM_L1L2XX_L3PHIC_dataarray_data_V_enb <= '1';
            else
              FM_L1L2XX_L3PHIC_dataarray_data_V_enb <= '0';
            end if;
            if (addr < (to_integer(unsigned(FM_L5L6XX_L3PHIC_nentries_V_dout(1))))) then -- Only read number of entries: Switch off in complete read out mode
              FM_L5L6XX_L3PHIC_dataarray_data_V_enb <= '1';
            else
              FM_L5L6XX_L3PHIC_dataarray_data_V_enb <= '0';
            end if;
          end if;
        end if;
        FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr <= std_logic_vector(to_unsigned(addr+(PAGE_OFFSET*(v_bx_cnt mod 2)),FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr'length));
        FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr <= std_logic_vector(to_unsigned(addr+(PAGE_OFFSET*(v_bx_cnt mod 2)),FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr'length));
        wait for 0 ns; -- Update signals
        -- Other writes ---------------------------------------
        if (addr >= MEM_READ_DELAY) then -- Take read dealy into account
          write(v_line, NOW, right, 20); -- NOW = current simulation time
          write(v_line, v_bx_cnt, right, 4);
          --write(v_line, string'("0x"), right, 4); hwrite(v_line, std_logic_vector(to_unsigned(addr,10)), right, 3);
          write(v_line, string'("0b"), right, 5);   write(v_line, reset, right, 1);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, FM_L1L2XX_L3PHIC_nentries_V_dout(0), right, 2);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, FM_L1L2XX_L3PHIC_nentries_V_dout(1), right, 2);
          write(v_line, string'("0b"), right, 3);   write(v_line, v_FM_L1L2XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-1), right, 1);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, std_logic_vector(unsigned(FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr)-to_unsigned(MEM_READ_DELAY,FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr'length)), right, 2);
          if (v_FM_L1L2XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-1)='1') then -- Only write if enable (delayed): Switch off in complete read out mode
            write(v_line, string'("0x"), right, 27); hwrite(v_line, FM_L1L2XX_L3PHIC_dataarray_data_V_dout, right, 12);
          else
            write(v_line, string'("0x"), right, 27);  write(v_line, string'("000000000000"), right, 12);
          end if;
          write(v_line, string'("0b"), right, 8);   write(v_line, MC_done, right, 1);
          write(v_line, string'("0b"), right, 13);  write(v_line, MC_bx_out_vld, right, 1);
          write(v_line, string'("0x"), right, 9);  hwrite(v_line, MC_bx_out, right, 1);
          writeline (file_out_L1L2, v_line); -- Write line
          write(v_line, NOW, right, 20); -- NOW = current simulation time
          write(v_line, v_bx_cnt, right, 4);
          --write(v_line, string'("0x"), right, 4); hwrite(v_line, std_logic_vector(to_unsigned(addr,10)), right, 3);
          write(v_line, string'("0b"), right, 5);   write(v_line, reset, right, 1);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, FM_L5L6XX_L3PHIC_nentries_V_dout(0), right, 2);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, FM_L5L6XX_L3PHIC_nentries_V_dout(1), right, 2);
          write(v_line, string'("0b"), right, 3);   write(v_line, v_FM_L5L6XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-1), right, 1);
          write(v_line, string'("0x"), right, 7);  hwrite(v_line, std_logic_vector(unsigned(FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr)-to_unsigned(MEM_READ_DELAY,FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr'length)), right, 2);
          if (v_FM_L5L6XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-1)='1') then -- Only write if enable (delayed): Switch off in complete read out mode
            write(v_line, string'("0x"), right, 27); hwrite(v_line, FM_L5L6XX_L3PHIC_dataarray_data_V_dout, right, 12);
          else
            write(v_line, string'("0x"), right, 27);  write(v_line, string'("000000000000"), right, 12);
          end if;
          write(v_line, string'("0b"), right, 8);   write(v_line, MC_done, right, 1);
          write(v_line, string'("0b"), right, 13);  write(v_line, MC_bx_out_vld, right, 1);
          write(v_line, string'("0x"), right, 9);  hwrite(v_line, MC_bx_out, right, 1);
          writeline (file_out_L5L6, v_line); -- Write line
        end if;
        v_FM_L1L2XX_L3PHIC_dataarray_data_V_enb_d :=  v_FM_L1L2XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-2 downto 0) & FM_L1L2XX_L3PHIC_dataarray_data_V_enb; -- Required delay
        v_FM_L5L6XX_L3PHIC_dataarray_data_V_enb_d :=  v_FM_L5L6XX_L3PHIC_dataarray_data_V_enb_d(MEM_READ_DELAY-2 downto 0) & FM_L5L6XX_L3PHIC_dataarray_data_V_enb; -- Required delay
        if (DEBUG=true and v_bx_cnt<=5 and addr<=10) then write(v_line, string'("v_bx_cnt: ")); write(v_line, v_bx_cnt); write(v_line, string'("   FM_L1L2XX_L3PHIC readaddr: ")); hwrite(v_line, FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr); write(v_line, string'(", dout: ")); hwrite(v_line, FM_L1L2XX_L3PHIC_dataarray_data_V_dout); writeline(output, v_line); end if;
        wait for CLK_PERIOD; -- Main time control
      end loop l_addr;
    end loop l_BX;
    file_close(file_out_L1L2);
    file_close(file_out_L5L6);
    assert false report "Simulation finished!" severity FAILURE;
  end process write_result;

  -- ########################### Instantiation ###########################
  -- Instantiate the Unit Under Test (UUT)
  i_top_tf : if INST_TOP_TF = 1 generate
    uut : entity work.top_tf
      port map(
        clk       => clk,
        reset     => reset,
        PR_start  => PR_start,
        PR_idle   => PR_idle,
        PR_ready  => PR_ready,
        PR_bx_in  => PR_bx_in,
        -- TrackletProjections input
        TPROJ_L3PHIC_dataarray_data_V_wea       => TPROJ_L3PHIC_dataarray_data_V_wea,
        TPROJ_L3PHIC_dataarray_data_V_writeaddr => TPROJ_L3PHIC_dataarray_data_V_writeaddr,
        TPROJ_L3PHIC_dataarray_data_V_din       => TPROJ_L3PHIC_dataarray_data_V_din,
        TPROJ_L3PHIC_nentries_V_we  => TPROJ_L3PHIC_nentries_V_we,
        TPROJ_L3PHIC_nentries_V_din => TPROJ_L3PHIC_nentries_V_din,
        -- VMStubsME input
        VMSME_L3PHIC17to24n1_dataarray_data_V_wea       => VMSME_L3PHIC17to24n1_dataarray_data_V_wea,
        VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr,
        VMSME_L3PHIC17to24n1_dataarray_data_V_din       => VMSME_L3PHIC17to24n1_dataarray_data_V_din,
        VMSME_L3PHIC17to24n1_nentries_V_we  => VMSME_L3PHIC17to24n1_nentries_V_we,
        VMSME_L3PHIC17to24n1_nentries_V_din => VMSME_L3PHIC17to24n1_nentries_V_din,
        -- AllStubs input
        AS_L3PHICn4_dataarray_data_V_wea       => AS_L3PHICn4_dataarray_data_V_wea,
        AS_L3PHICn4_dataarray_data_V_writeaddr => AS_L3PHICn4_dataarray_data_V_writeaddr,
        AS_L3PHICn4_dataarray_data_V_din       => AS_L3PHICn4_dataarray_data_V_din,
        AS_L3PHICn4_nentries_V_we  => AS_L3PHICn4_nentries_V_we,
        AS_L3PHICn4_nentries_V_din => AS_L3PHICn4_nentries_V_din,
        -- FullMatches output
        FM_L1L2XX_L3PHIC_dataarray_data_V_enb      => FM_L1L2XX_L3PHIC_dataarray_data_V_enb,
        FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr => FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L1L2XX_L3PHIC_dataarray_data_V_dout     => FM_L1L2XX_L3PHIC_dataarray_data_V_dout,
        FM_L1L2XX_L3PHIC_nentries_V_dout            => FM_L1L2XX_L3PHIC_nentries_V_dout,
        FM_L5L6XX_L3PHIC_dataarray_data_V_enb      => FM_L5L6XX_L3PHIC_dataarray_data_V_enb,
        FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr => FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L5L6XX_L3PHIC_dataarray_data_V_dout     => FM_L5L6XX_L3PHIC_dataarray_data_V_dout,
        FM_L5L6XX_L3PHIC_nentries_V_dout            => FM_L5L6XX_L3PHIC_nentries_V_dout,
        -- MatchCalculator output
        MC_bx_out     => MC_bx_out,
        MC_bx_out_vld => MC_bx_out_vld,
        MC_done       => MC_done );
  end generate;

  i_top_tf_full : if INST_TOP_TF = 2 generate
    uut : entity work.top_tf_full
      port map(
        clk       => clk,
        reset     => reset,
        PR_start  => PR_start,
        PR_idle   => PR_idle,
        PR_ready  => PR_ready,
        PR_bx_in  => PR_bx_in,
        -- TrackletProjections input
        TPROJ_L3PHIC_dataarray_data_V_wea       => TPROJ_L3PHIC_dataarray_data_V_wea,
        TPROJ_L3PHIC_dataarray_data_V_writeaddr => TPROJ_L3PHIC_dataarray_data_V_writeaddr,
        TPROJ_L3PHIC_dataarray_data_V_din       => TPROJ_L3PHIC_dataarray_data_V_din,
        TPROJ_L3PHIC_nentries_V_we  => TPROJ_L3PHIC_nentries_V_we,
        TPROJ_L3PHIC_nentries_V_din => TPROJ_L3PHIC_nentries_V_din,
        -- VMStubsME input
        VMSME_L3PHIC17to24n1_dataarray_data_V_wea       => VMSME_L3PHIC17to24n1_dataarray_data_V_wea,
        VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr,
        VMSME_L3PHIC17to24n1_dataarray_data_V_din       => VMSME_L3PHIC17to24n1_dataarray_data_V_din,
        VMSME_L3PHIC17to24n1_nentries_V_we  => VMSME_L3PHIC17to24n1_nentries_V_we,
        VMSME_L3PHIC17to24n1_nentries_V_din => VMSME_L3PHIC17to24n1_nentries_V_din,
        -- AllStubs input
        AS_L3PHICn4_dataarray_data_V_wea       => AS_L3PHICn4_dataarray_data_V_wea,
        AS_L3PHICn4_dataarray_data_V_writeaddr => AS_L3PHICn4_dataarray_data_V_writeaddr,
        AS_L3PHICn4_dataarray_data_V_din       => AS_L3PHICn4_dataarray_data_V_din,
        AS_L3PHICn4_nentries_V_we  => AS_L3PHICn4_nentries_V_we,
        AS_L3PHICn4_nentries_V_din => AS_L3PHICn4_nentries_V_din,
        -- VMProjection output
        VMPROJ_L3PHIC17to24_dataarray_data_V_wea       => VMPROJ_L3PHIC17to24_dataarray_data_V_wea,
        VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr => VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr,
        VMPROJ_L3PHIC17to24_dataarray_data_V_din       => VMPROJ_L3PHIC17to24_dataarray_data_V_din,
        --VMPROJ_L3PHIC17to24_nentries_V_we              => VMPROJ_L3PHIC17to24_nentries_V_we,
        --VMPROJ_L3PHIC17to24_nentries_V_din             => VMPROJ_L3PHIC17to24_nentries_V_din,
        -- AllProjection output
        AP_L3PHIC_dataarray_data_V_wea       => AP_L3PHIC_dataarray_data_V_wea,
        AP_L3PHIC_dataarray_data_V_writeaddr => AP_L3PHIC_dataarray_data_V_writeaddr,
        AP_L3PHIC_dataarray_data_V_din       => AP_L3PHIC_dataarray_data_V_din,
        --AP_L3PHIC_nentries_V_we              => AP_L3PHIC_nentries_V_we,
        --AP_L3PHIC_nentries_V_din             => AP_L3PHIC_nentries_V_din,
        -- ProjectionRouter output
        PR_bx_out     => PR_bx_out,
        PR_bx_out_vld => PR_bx_out_vld,
        PR_done       => PR_done,
        -- CandidateMatch output
        CM_L3PHIC17to24_dataarray_data_V_wea       => CM_L3PHIC17to24_dataarray_data_V_wea,
        CM_L3PHIC17to24_dataarray_data_V_writeaddr => CM_L3PHIC17to24_dataarray_data_V_writeaddr,
        CM_L3PHIC17to24_dataarray_data_V_din       => CM_L3PHIC17to24_dataarray_data_V_din,
        --CM_L3PHIC17to24_nentries_V_we              => CM_L3PHIC17to24_nentries_V_we,
        --CM_L3PHIC17to24_nentries_V_din             => CM_L3PHIC17to24_nentries_V_din,
        -- MatchEngine output
        ME_bx_out     => ME_bx_out,
        ME_bx_out_vld => ME_bx_out_vld,
        ME_all_done   => ME_all_done,
        -- FullMatches output
        FM_L1L2XX_L3PHIC_dataarray_data_V_enb      => FM_L1L2XX_L3PHIC_dataarray_data_V_enb,
        FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr => FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L1L2XX_L3PHIC_dataarray_data_V_dout     => FM_L1L2XX_L3PHIC_dataarray_data_V_dout,
        FM_L1L2XX_L3PHIC_nentries_V_dout           => FM_L1L2XX_L3PHIC_nentries_V_dout,
        FM_L5L6XX_L3PHIC_dataarray_data_V_enb      => FM_L5L6XX_L3PHIC_dataarray_data_V_enb,
        FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr => FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L5L6XX_L3PHIC_dataarray_data_V_dout     => FM_L5L6XX_L3PHIC_dataarray_data_V_dout,
        FM_L5L6XX_L3PHIC_nentries_V_dout           => FM_L5L6XX_L3PHIC_nentries_V_dout,
        -- MatchCalculator output
        MC_bx_out     => MC_bx_out,
        MC_bx_out_vld => MC_bx_out_vld,
        MC_done       => MC_done );
    --! @brief TextIO process for writting the output ---------------------------------------
    write_result_AP : process
      variable v_bx_cnt      : integer       := -1; --! BX counter
    begin
      wait until PR_start = '1'; -- Wait to start
      write_header_line(FILE_OUT_AP, "AP_L3PHIC_dataarray_data_V_din", 8);
      l_BX : while v_bx_cnt <= MAX_EVENTS-1 loop
        if (AP_L3PHIC_dataarray_data_V_writeaddr(6 downto 0) = b"000_0000") and
           (AP_L3PHIC_dataarray_data_V_wea = '1') then -- Start new event assuming all addr behave the same
          v_bx_cnt := v_bx_cnt + 1;
        end if;
        if (AP_L3PHIC_dataarray_data_V_wea='1') then -- Only write valid data
                --or AP_L3PHIC_nentries_V_we(0)='1' or AP_L3PHIC_nentries_V_we(1)='1' or
                --AP_L3PHIC_nentries_V_we(2)='1' or AP_L3PHIC_nentries_V_we(3)='1' or AP_L3PHIC_nentries_V_we(4)='1' or
                --AP_L3PHIC_nentries_V_we(5)='1' or AP_L3PHIC_nentries_V_we(6)='1' or AP_L3PHIC_nentries_V_we(7)='1') then -- Only write valid data
          write_emData_line_8p(reset, v_bx_cnt, PR_done, PR_bx_out, PR_bx_out_vld, FILE_OUT_AP, "AP_L3PHIC_dataarray_data_V_din",
                               AP_L3PHIC_dataarray_data_V_din, AP_L3PHIC_dataarray_data_V_wea, AP_L3PHIC_dataarray_data_V_writeaddr,
                               (others => (others => '0')), (others => '0') );--AP_L3PHIC_nentries_V_din, AP_L3PHIC_nentries_V_we );
        end if;
        wait for CLK_PERIOD; -- Main time control
      end loop l_BX;
      wait;
    end process write_result_AP;
    --! @brief TextIO process for writting the output ---------------------------------------
    write_result_VMP : process
      variable v_bx_cnt      : integer       := -1; --! BX counter
      variable myarray2_8b   : t_myarray2_8b := (others => (others => '0')); -- Temporary array to avoid sim error
      variable myarray2_1b   : t_myarray2_1b := (others => '0'); -- Temporary array to avoid sim error
      variable v_addr_d1     : t_myarray8_8b := (others => (others => '0')); -- Delayed address
    begin
      wait until PR_start = '1'; -- Wait to start
      l_copies_header : for cp in 0 to N_ME_IN_CHAIN-1 loop -- 0 to 7
        write_header_line(FILE_OUT_VMP(cp), "VMPROJ_L3PHIC17to24_dataarray_data_V_din", 2);
      end loop l_copies_header;
      l_BX : while v_bx_cnt <= MAX_EVENTS-1 loop
        if (VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr(0)(6 downto 0) = b"000_0000") and
           v_addr_d1(0)(7) /= VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr(0)(7) then -- Start new event assuming all addr behave the same
          v_bx_cnt := v_bx_cnt + 1;
        end if;
        l_copies : for cp in 0 to N_ME_IN_CHAIN-1 loop -- 0 to 7
          if (VMPROJ_L3PHIC17to24_dataarray_data_V_wea(cp)='1') then -- Only write valid data
          --if (VMPROJ_L3PHIC17to24_dataarray_data_V_wea(cp)='1' or VMPROJ_L3PHIC17to24_nentries_V_we(0)(cp)='1' or VMPROJ_L3PHIC17to24_nentries_V_we(1)(cp)='1') then -- Only write valid data
            --myarray2_8b := (VMPROJ_L3PHIC17to24_nentries_V_din(0)(cp)) & (VMPROJ_L3PHIC17to24_nentries_V_din(1)(cp)); -- Needed to avoid sim error (casting does not work)
            --myarray2_1b := (VMPROJ_L3PHIC17to24_nentries_V_we(0)(cp))  & (VMPROJ_L3PHIC17to24_nentries_V_we(1)(cp));  -- Needed to avoid sim error (casting does not work)
            write_emData_line_2p(reset, v_bx_cnt, PR_done, PR_bx_out, PR_bx_out_vld, FILE_OUT_VMP(cp), "VMPROJ_L3PHIC17to24_dataarray_data_V_din",
                                 VMPROJ_L3PHIC17to24_dataarray_data_V_din(cp), VMPROJ_L3PHIC17to24_dataarray_data_V_wea(cp), VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr(cp),
                                 myarray2_8b, myarray2_1b );
          end if;
        end loop l_copies;
        v_addr_d1 := VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr; -- Delay the address
        wait for CLK_PERIOD; -- Main time control
      end loop l_BX;
      wait;
    end process write_result_VMP;
    --! @brief TextIO process for writting the output ---------------------------------------
    write_result_CM : process
      variable v_bx_cnt    : integer       := -1; --! BX counter
      variable myarray2_8b : t_myarray2_8b := (others => (others => '0')); -- Temporary array to avoid sim error
      variable myarray2_1b : t_myarray2_1b := (others => '0'); -- Temporary array to avoid sim error
      variable v_addr_d1   : t_myarray8_8b := (others => (others => '0')); -- Delayed address
    begin
      wait until PR_done = '1'; -- Wait to start = ME_start
      l_copies_header : for cp in 0 to N_ME_IN_CHAIN-1 loop -- 0 to 7
        write_header_line(FILE_OUT_CM(cp), "CM_L3PHIC17to24_dataarray_data_V_din", 2);
      end loop l_copies_header;
      l_BX : while v_bx_cnt <= MAX_EVENTS-1 loop
        if (CM_L3PHIC17to24_dataarray_data_V_writeaddr(0)(6 downto 0) = b"000_0000") and
           v_addr_d1(0)(7) /= CM_L3PHIC17to24_dataarray_data_V_writeaddr(0)(7) then -- Start new event assuming all addr behave the same
          v_bx_cnt := v_bx_cnt + 1;
        end if;
        l_copies : for cp in 0 to N_ME_IN_CHAIN-1 loop -- 0 to 7
          if (CM_L3PHIC17to24_dataarray_data_V_wea(cp)='1') then
          --if (CM_L3PHIC17to24_dataarray_data_V_wea(cp)='1' or CM_L3PHIC17to24_nentries_V_we(0)(cp)='1' or CM_L3PHIC17to24_nentries_V_we(1)(cp)='1') then -- Only write valid data
            --myarray2_8b := (CM_L3PHIC17to24_nentries_V_din(0)(cp)) & (CM_L3PHIC17to24_nentries_V_din(1)(cp)); -- Needed to avoid sim error (casting does not work)
            --myarray2_1b := (CM_L3PHIC17to24_nentries_V_we(0)(cp))  & (CM_L3PHIC17to24_nentries_V_we(1)(cp));  -- Needed to avoid sim error (casting does not work)
            write_emData_line_2p(reset, v_bx_cnt, ME_all_done, ME_bx_out(cp), ME_bx_out_vld(cp), FILE_OUT_CM(cp), "CM_L3PHIC17to24_dataarray_data_V_din",
                                 CM_L3PHIC17to24_dataarray_data_V_din(cp), CM_L3PHIC17to24_dataarray_data_V_wea(cp), CM_L3PHIC17to24_dataarray_data_V_writeaddr(cp),
                                 myarray2_8b, myarray2_1b );
          end if;
        end loop l_copies;
        v_addr_d1 := CM_L3PHIC17to24_dataarray_data_V_writeaddr; -- Delay the address
        wait for CLK_PERIOD; -- Main time control
      end loop l_BX;
      wait;
    end process write_result_CM;
  end generate;

  i_others : if INST_TOP_TF = 0 generate
    uut : entity work.SectorProcessor
      port map(
        clk        => clk,
        reset      => reset,
        en_proc                => PR_start,
        bx_in_ProjectionRouter => PR_bx_in,
        bx_out_MatchCalculator     => MC_bx_out,
        bx_out_MatchCalculator_vld => MC_bx_out_vld,
        MatchCalculator_done       => MC_done,
        TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(0),
        TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(0),
        TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(0),
        TPROJ_L1L2XXF_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(0),
        TPROJ_L1L2XXF_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(0),
        TPROJ_L1L2XXF_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(0),
        TPROJ_L1L2XXF_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(0),
        TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(1),
        TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(1),
        TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(1),
        TPROJ_L1L2XXG_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(1),
        TPROJ_L1L2XXG_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(1),
        TPROJ_L1L2XXG_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(1),
        TPROJ_L1L2XXG_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(1),
        TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(2),
        TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(2),
        TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(2),
        TPROJ_L1L2XXH_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(2),
        TPROJ_L1L2XXH_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(2),
        TPROJ_L1L2XXH_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(2),
        TPROJ_L1L2XXH_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(2),
        TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(3),
        TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(3),
        TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(3),
        TPROJ_L1L2XXI_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(3),
        TPROJ_L1L2XXI_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(3),
        TPROJ_L1L2XXI_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(3),
        TPROJ_L1L2XXI_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(3),
        TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(4),
        TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(4),
        TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(4),
        TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(4),
        TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(4),
        TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(4),
        TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(4),
        TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(5),
        TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(5),
        TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(5),
        TPROJ_L5L6XXB_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(5),
        TPROJ_L5L6XXB_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(5),
        TPROJ_L5L6XXB_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(5),
        TPROJ_L5L6XXB_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(5),
        TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(6),
        TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(6),
        TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(6),
        TPROJ_L5L6XXC_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(6),
        TPROJ_L5L6XXC_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(6),
        TPROJ_L5L6XXC_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(6),
        TPROJ_L5L6XXC_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(6),
        TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_wea       =>           TPROJ_L3PHIC_dataarray_data_V_wea(7),
        TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_writeaddr =>     TPROJ_L3PHIC_dataarray_data_V_writeaddr(7),
        TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_din       =>           TPROJ_L3PHIC_dataarray_data_V_din(7),
        TPROJ_L5L6XXD_L3PHIC_nentries_0_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(0)(7),
        TPROJ_L5L6XXD_L3PHIC_nentries_0_V_din =>                        TPROJ_L3PHIC_nentries_V_din(0)(7),
        TPROJ_L5L6XXD_L3PHIC_nentries_1_V_we  =>                         TPROJ_L3PHIC_nentries_V_we(1)(7),
        TPROJ_L5L6XXD_L3PHIC_nentries_1_V_din =>                        TPROJ_L3PHIC_nentries_V_din(1)(7),
        VMSME_L3PHIC17n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(0),
        VMSME_L3PHIC17n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(0),
        VMSME_L3PHIC17n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(0),
        VMSME_L3PHIC17n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(0),
        VMSME_L3PHIC17n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(0),
        VMSME_L3PHIC17n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(0),
        VMSME_L3PHIC17n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(0),
        VMSME_L3PHIC17n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(0),
        VMSME_L3PHIC17n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(0),
        VMSME_L3PHIC17n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(0),
        VMSME_L3PHIC17n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(0),
        VMSME_L3PHIC17n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(0),
        VMSME_L3PHIC17n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(0),
        VMSME_L3PHIC17n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(0),
        VMSME_L3PHIC17n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(0),
        VMSME_L3PHIC17n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(0),
        VMSME_L3PHIC17n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(0),
        VMSME_L3PHIC17n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(0),
        VMSME_L3PHIC17n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(0),
        VMSME_L3PHIC17n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(0),
        VMSME_L3PHIC17n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(0),
        VMSME_L3PHIC17n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(0),
        VMSME_L3PHIC17n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(0),
        VMSME_L3PHIC17n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(0),
        VMSME_L3PHIC17n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(0),
        VMSME_L3PHIC17n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(0),
        VMSME_L3PHIC17n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(0),
        VMSME_L3PHIC17n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(0),
        VMSME_L3PHIC17n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(0),
        VMSME_L3PHIC17n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(0),
        VMSME_L3PHIC17n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(0),
        VMSME_L3PHIC17n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(0),
        VMSME_L3PHIC17n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(0),
        VMSME_L3PHIC17n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(0),
        VMSME_L3PHIC17n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(0),
        VMSME_L3PHIC17n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(0),
        VMSME_L3PHIC17n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(0),
        VMSME_L3PHIC17n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(0),
        VMSME_L3PHIC17n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(0),
        VMSME_L3PHIC17n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(0),
        VMSME_L3PHIC17n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(0),
        VMSME_L3PHIC17n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(0),
        VMSME_L3PHIC17n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(0),
        VMSME_L3PHIC17n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(0),
        VMSME_L3PHIC17n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(0),
        VMSME_L3PHIC17n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(0),
        VMSME_L3PHIC17n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(0),
        VMSME_L3PHIC17n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(0),
        VMSME_L3PHIC17n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(0),
        VMSME_L3PHIC17n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(0),
        VMSME_L3PHIC17n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(0),
        VMSME_L3PHIC17n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(0),
        VMSME_L3PHIC17n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(0),
        VMSME_L3PHIC17n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(0),
        VMSME_L3PHIC17n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(0),
        VMSME_L3PHIC17n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(0),
        VMSME_L3PHIC17n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(0),
        VMSME_L3PHIC17n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(0),
        VMSME_L3PHIC17n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(0),
        VMSME_L3PHIC17n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(0),
        VMSME_L3PHIC17n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(0),
        VMSME_L3PHIC17n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(0),
        VMSME_L3PHIC17n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(0),
        VMSME_L3PHIC17n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(0),
        VMSME_L3PHIC17n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(0),
        VMSME_L3PHIC17n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(0),
        VMSME_L3PHIC17n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(0),
        VMSME_L3PHIC17n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(0),
        VMSME_L3PHIC17n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(0),
        VMSME_L3PHIC17n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(0),
        VMSME_L3PHIC17n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(0),
        VMSME_L3PHIC17n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(0),
        VMSME_L3PHIC17n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(0),
        VMSME_L3PHIC17n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(0),
        VMSME_L3PHIC17n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(0),
        VMSME_L3PHIC17n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(0),
        VMSME_L3PHIC17n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(0),
        VMSME_L3PHIC17n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(0),
        VMSME_L3PHIC17n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(0),
        VMSME_L3PHIC17n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(0),
        VMSME_L3PHIC17n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(0),
        VMSME_L3PHIC17n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(0),
        VMSME_L3PHIC17n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(0),
        VMSME_L3PHIC17n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(0),
        VMSME_L3PHIC17n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(0),
        VMSME_L3PHIC17n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(0),
        VMSME_L3PHIC17n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(0),
        VMSME_L3PHIC17n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(0),
        VMSME_L3PHIC17n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(0),
        VMSME_L3PHIC17n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(0),
        VMSME_L3PHIC17n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(0),
        VMSME_L3PHIC17n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(0),
        VMSME_L3PHIC17n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(0),
        VMSME_L3PHIC17n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(0),
        VMSME_L3PHIC17n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(0),
        VMSME_L3PHIC17n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(0),
        VMSME_L3PHIC17n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(0),
        VMSME_L3PHIC17n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(0),
        VMSME_L3PHIC17n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(0),
        VMSME_L3PHIC17n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(0),
        VMSME_L3PHIC17n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(0),
        VMSME_L3PHIC17n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(0),
        VMSME_L3PHIC17n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(0),
        VMSME_L3PHIC17n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(0),
        VMSME_L3PHIC17n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(0),
        VMSME_L3PHIC17n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(0),
        VMSME_L3PHIC17n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(0),
        VMSME_L3PHIC17n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(0),
        VMSME_L3PHIC17n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(0),
        VMSME_L3PHIC17n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(0),
        VMSME_L3PHIC17n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(0),
        VMSME_L3PHIC17n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(0),
        VMSME_L3PHIC17n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(0),
        VMSME_L3PHIC17n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(0),
        VMSME_L3PHIC17n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(0),
        VMSME_L3PHIC17n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(0),
        VMSME_L3PHIC17n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(0),
        VMSME_L3PHIC17n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(0),
        VMSME_L3PHIC17n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(0),
        VMSME_L3PHIC17n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(0),
        VMSME_L3PHIC17n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(0),
        VMSME_L3PHIC17n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(0),
        VMSME_L3PHIC17n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(0),
        VMSME_L3PHIC17n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(0),
        VMSME_L3PHIC17n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(0),
        VMSME_L3PHIC17n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(0),
        VMSME_L3PHIC17n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(0),
        VMSME_L3PHIC17n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(0),
        VMSME_L3PHIC17n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(0),
        VMSME_L3PHIC17n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(0),
        VMSME_L3PHIC17n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(0),
        VMSME_L3PHIC18n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(1),
        VMSME_L3PHIC18n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(1),
        VMSME_L3PHIC18n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(1),
        VMSME_L3PHIC18n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(1),
        VMSME_L3PHIC18n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(1),
        VMSME_L3PHIC18n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(1),
        VMSME_L3PHIC18n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(1),
        VMSME_L3PHIC18n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(1),
        VMSME_L3PHIC18n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(1),
        VMSME_L3PHIC18n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(1),
        VMSME_L3PHIC18n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(1),
        VMSME_L3PHIC18n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(1),
        VMSME_L3PHIC18n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(1),
        VMSME_L3PHIC18n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(1),
        VMSME_L3PHIC18n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(1),
        VMSME_L3PHIC18n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(1),
        VMSME_L3PHIC18n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(1),
        VMSME_L3PHIC18n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(1),
        VMSME_L3PHIC18n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(1),
        VMSME_L3PHIC18n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(1),
        VMSME_L3PHIC18n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(1),
        VMSME_L3PHIC18n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(1),
        VMSME_L3PHIC18n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(1),
        VMSME_L3PHIC18n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(1),
        VMSME_L3PHIC18n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(1),
        VMSME_L3PHIC18n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(1),
        VMSME_L3PHIC18n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(1),
        VMSME_L3PHIC18n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(1),
        VMSME_L3PHIC18n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(1),
        VMSME_L3PHIC18n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(1),
        VMSME_L3PHIC18n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(1),
        VMSME_L3PHIC18n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(1),
        VMSME_L3PHIC18n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(1),
        VMSME_L3PHIC18n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(1),
        VMSME_L3PHIC18n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(1),
        VMSME_L3PHIC18n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(1),
        VMSME_L3PHIC18n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(1),
        VMSME_L3PHIC18n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(1),
        VMSME_L3PHIC18n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(1),
        VMSME_L3PHIC18n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(1),
        VMSME_L3PHIC18n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(1),
        VMSME_L3PHIC18n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(1),
        VMSME_L3PHIC18n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(1),
        VMSME_L3PHIC18n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(1),
        VMSME_L3PHIC18n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(1),
        VMSME_L3PHIC18n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(1),
        VMSME_L3PHIC18n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(1),
        VMSME_L3PHIC18n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(1),
        VMSME_L3PHIC18n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(1),
        VMSME_L3PHIC18n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(1),
        VMSME_L3PHIC18n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(1),
        VMSME_L3PHIC18n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(1),
        VMSME_L3PHIC18n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(1),
        VMSME_L3PHIC18n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(1),
        VMSME_L3PHIC18n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(1),
        VMSME_L3PHIC18n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(1),
        VMSME_L3PHIC18n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(1),
        VMSME_L3PHIC18n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(1),
        VMSME_L3PHIC18n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(1),
        VMSME_L3PHIC18n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(1),
        VMSME_L3PHIC18n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(1),
        VMSME_L3PHIC18n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(1),
        VMSME_L3PHIC18n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(1),
        VMSME_L3PHIC18n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(1),
        VMSME_L3PHIC18n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(1),
        VMSME_L3PHIC18n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(1),
        VMSME_L3PHIC18n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(1),
        VMSME_L3PHIC18n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(1),
        VMSME_L3PHIC18n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(1),
        VMSME_L3PHIC18n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(1),
        VMSME_L3PHIC18n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(1),
        VMSME_L3PHIC18n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(1),
        VMSME_L3PHIC18n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(1),
        VMSME_L3PHIC18n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(1),
        VMSME_L3PHIC18n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(1),
        VMSME_L3PHIC18n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(1),
        VMSME_L3PHIC18n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(1),
        VMSME_L3PHIC18n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(1),
        VMSME_L3PHIC18n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(1),
        VMSME_L3PHIC18n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(1),
        VMSME_L3PHIC18n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(1),
        VMSME_L3PHIC18n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(1),
        VMSME_L3PHIC18n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(1),
        VMSME_L3PHIC18n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(1),
        VMSME_L3PHIC18n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(1),
        VMSME_L3PHIC18n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(1),
        VMSME_L3PHIC18n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(1),
        VMSME_L3PHIC18n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(1),
        VMSME_L3PHIC18n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(1),
        VMSME_L3PHIC18n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(1),
        VMSME_L3PHIC18n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(1),
        VMSME_L3PHIC18n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(1),
        VMSME_L3PHIC18n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(1),
        VMSME_L3PHIC18n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(1),
        VMSME_L3PHIC18n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(1),
        VMSME_L3PHIC18n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(1),
        VMSME_L3PHIC18n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(1),
        VMSME_L3PHIC18n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(1),
        VMSME_L3PHIC18n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(1),
        VMSME_L3PHIC18n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(1),
        VMSME_L3PHIC18n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(1),
        VMSME_L3PHIC18n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(1),
        VMSME_L3PHIC18n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(1),
        VMSME_L3PHIC18n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(1),
        VMSME_L3PHIC18n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(1),
        VMSME_L3PHIC18n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(1),
        VMSME_L3PHIC18n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(1),
        VMSME_L3PHIC18n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(1),
        VMSME_L3PHIC18n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(1),
        VMSME_L3PHIC18n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(1),
        VMSME_L3PHIC18n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(1),
        VMSME_L3PHIC18n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(1),
        VMSME_L3PHIC18n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(1),
        VMSME_L3PHIC18n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(1),
        VMSME_L3PHIC18n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(1),
        VMSME_L3PHIC18n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(1),
        VMSME_L3PHIC18n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(1),
        VMSME_L3PHIC18n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(1),
        VMSME_L3PHIC18n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(1),
        VMSME_L3PHIC18n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(1),
        VMSME_L3PHIC18n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(1),
        VMSME_L3PHIC18n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(1),
        VMSME_L3PHIC18n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(1),
        VMSME_L3PHIC18n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(1),
        VMSME_L3PHIC18n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(1),
        VMSME_L3PHIC18n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(1),
        VMSME_L3PHIC18n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(1),
        VMSME_L3PHIC18n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(1),
        VMSME_L3PHIC18n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(1),
        VMSME_L3PHIC18n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(1),
        VMSME_L3PHIC18n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(1),
        VMSME_L3PHIC19n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(2),
        VMSME_L3PHIC19n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(2),
        VMSME_L3PHIC19n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(2),
        VMSME_L3PHIC19n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(2),
        VMSME_L3PHIC19n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(2),
        VMSME_L3PHIC19n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(2),
        VMSME_L3PHIC19n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(2),
        VMSME_L3PHIC19n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(2),
        VMSME_L3PHIC19n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(2),
        VMSME_L3PHIC19n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(2),
        VMSME_L3PHIC19n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(2),
        VMSME_L3PHIC19n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(2),
        VMSME_L3PHIC19n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(2),
        VMSME_L3PHIC19n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(2),
        VMSME_L3PHIC19n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(2),
        VMSME_L3PHIC19n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(2),
        VMSME_L3PHIC19n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(2),
        VMSME_L3PHIC19n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(2),
        VMSME_L3PHIC19n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(2),
        VMSME_L3PHIC19n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(2),
        VMSME_L3PHIC19n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(2),
        VMSME_L3PHIC19n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(2),
        VMSME_L3PHIC19n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(2),
        VMSME_L3PHIC19n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(2),
        VMSME_L3PHIC19n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(2),
        VMSME_L3PHIC19n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(2),
        VMSME_L3PHIC19n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(2),
        VMSME_L3PHIC19n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(2),
        VMSME_L3PHIC19n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(2),
        VMSME_L3PHIC19n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(2),
        VMSME_L3PHIC19n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(2),
        VMSME_L3PHIC19n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(2),
        VMSME_L3PHIC19n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(2),
        VMSME_L3PHIC19n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(2),
        VMSME_L3PHIC19n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(2),
        VMSME_L3PHIC19n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(2),
        VMSME_L3PHIC19n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(2),
        VMSME_L3PHIC19n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(2),
        VMSME_L3PHIC19n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(2),
        VMSME_L3PHIC19n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(2),
        VMSME_L3PHIC19n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(2),
        VMSME_L3PHIC19n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(2),
        VMSME_L3PHIC19n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(2),
        VMSME_L3PHIC19n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(2),
        VMSME_L3PHIC19n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(2),
        VMSME_L3PHIC19n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(2),
        VMSME_L3PHIC19n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(2),
        VMSME_L3PHIC19n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(2),
        VMSME_L3PHIC19n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(2),
        VMSME_L3PHIC19n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(2),
        VMSME_L3PHIC19n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(2),
        VMSME_L3PHIC19n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(2),
        VMSME_L3PHIC19n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(2),
        VMSME_L3PHIC19n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(2),
        VMSME_L3PHIC19n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(2),
        VMSME_L3PHIC19n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(2),
        VMSME_L3PHIC19n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(2),
        VMSME_L3PHIC19n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(2),
        VMSME_L3PHIC19n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(2),
        VMSME_L3PHIC19n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(2),
        VMSME_L3PHIC19n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(2),
        VMSME_L3PHIC19n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(2),
        VMSME_L3PHIC19n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(2),
        VMSME_L3PHIC19n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(2),
        VMSME_L3PHIC19n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(2),
        VMSME_L3PHIC19n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(2),
        VMSME_L3PHIC19n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(2),
        VMSME_L3PHIC19n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(2),
        VMSME_L3PHIC19n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(2),
        VMSME_L3PHIC19n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(2),
        VMSME_L3PHIC19n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(2),
        VMSME_L3PHIC19n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(2),
        VMSME_L3PHIC19n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(2),
        VMSME_L3PHIC19n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(2),
        VMSME_L3PHIC19n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(2),
        VMSME_L3PHIC19n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(2),
        VMSME_L3PHIC19n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(2),
        VMSME_L3PHIC19n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(2),
        VMSME_L3PHIC19n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(2),
        VMSME_L3PHIC19n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(2),
        VMSME_L3PHIC19n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(2),
        VMSME_L3PHIC19n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(2),
        VMSME_L3PHIC19n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(2),
        VMSME_L3PHIC19n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(2),
        VMSME_L3PHIC19n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(2),
        VMSME_L3PHIC19n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(2),
        VMSME_L3PHIC19n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(2),
        VMSME_L3PHIC19n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(2),
        VMSME_L3PHIC19n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(2),
        VMSME_L3PHIC19n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(2),
        VMSME_L3PHIC19n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(2),
        VMSME_L3PHIC19n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(2),
        VMSME_L3PHIC19n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(2),
        VMSME_L3PHIC19n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(2),
        VMSME_L3PHIC19n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(2),
        VMSME_L3PHIC19n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(2),
        VMSME_L3PHIC19n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(2),
        VMSME_L3PHIC19n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(2),
        VMSME_L3PHIC19n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(2),
        VMSME_L3PHIC19n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(2),
        VMSME_L3PHIC19n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(2),
        VMSME_L3PHIC19n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(2),
        VMSME_L3PHIC19n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(2),
        VMSME_L3PHIC19n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(2),
        VMSME_L3PHIC19n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(2),
        VMSME_L3PHIC19n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(2),
        VMSME_L3PHIC19n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(2),
        VMSME_L3PHIC19n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(2),
        VMSME_L3PHIC19n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(2),
        VMSME_L3PHIC19n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(2),
        VMSME_L3PHIC19n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(2),
        VMSME_L3PHIC19n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(2),
        VMSME_L3PHIC19n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(2),
        VMSME_L3PHIC19n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(2),
        VMSME_L3PHIC19n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(2),
        VMSME_L3PHIC19n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(2),
        VMSME_L3PHIC19n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(2),
        VMSME_L3PHIC19n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(2),
        VMSME_L3PHIC19n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(2),
        VMSME_L3PHIC19n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(2),
        VMSME_L3PHIC19n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(2),
        VMSME_L3PHIC19n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(2),
        VMSME_L3PHIC19n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(2),
        VMSME_L3PHIC19n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(2),
        VMSME_L3PHIC19n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(2),
        VMSME_L3PHIC19n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(2),
        VMSME_L3PHIC19n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(2),
        VMSME_L3PHIC19n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(2),
        VMSME_L3PHIC19n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(2),
        VMSME_L3PHIC19n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(2),
        VMSME_L3PHIC19n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(2),
        VMSME_L3PHIC20n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(3),
        VMSME_L3PHIC20n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(3),
        VMSME_L3PHIC20n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(3),
        VMSME_L3PHIC20n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(3),
        VMSME_L3PHIC20n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(3),
        VMSME_L3PHIC20n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(3),
        VMSME_L3PHIC20n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(3),
        VMSME_L3PHIC20n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(3),
        VMSME_L3PHIC20n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(3),
        VMSME_L3PHIC20n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(3),
        VMSME_L3PHIC20n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(3),
        VMSME_L3PHIC20n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(3),
        VMSME_L3PHIC20n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(3),
        VMSME_L3PHIC20n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(3),
        VMSME_L3PHIC20n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(3),
        VMSME_L3PHIC20n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(3),
        VMSME_L3PHIC20n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(3),
        VMSME_L3PHIC20n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(3),
        VMSME_L3PHIC20n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(3),
        VMSME_L3PHIC20n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(3),
        VMSME_L3PHIC20n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(3),
        VMSME_L3PHIC20n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(3),
        VMSME_L3PHIC20n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(3),
        VMSME_L3PHIC20n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(3),
        VMSME_L3PHIC20n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(3),
        VMSME_L3PHIC20n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(3),
        VMSME_L3PHIC20n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(3),
        VMSME_L3PHIC20n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(3),
        VMSME_L3PHIC20n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(3),
        VMSME_L3PHIC20n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(3),
        VMSME_L3PHIC20n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(3),
        VMSME_L3PHIC20n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(3),
        VMSME_L3PHIC20n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(3),
        VMSME_L3PHIC20n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(3),
        VMSME_L3PHIC20n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(3),
        VMSME_L3PHIC20n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(3),
        VMSME_L3PHIC20n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(3),
        VMSME_L3PHIC20n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(3),
        VMSME_L3PHIC20n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(3),
        VMSME_L3PHIC20n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(3),
        VMSME_L3PHIC20n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(3),
        VMSME_L3PHIC20n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(3),
        VMSME_L3PHIC20n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(3),
        VMSME_L3PHIC20n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(3),
        VMSME_L3PHIC20n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(3),
        VMSME_L3PHIC20n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(3),
        VMSME_L3PHIC20n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(3),
        VMSME_L3PHIC20n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(3),
        VMSME_L3PHIC20n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(3),
        VMSME_L3PHIC20n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(3),
        VMSME_L3PHIC20n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(3),
        VMSME_L3PHIC20n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(3),
        VMSME_L3PHIC20n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(3),
        VMSME_L3PHIC20n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(3),
        VMSME_L3PHIC20n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(3),
        VMSME_L3PHIC20n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(3),
        VMSME_L3PHIC20n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(3),
        VMSME_L3PHIC20n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(3),
        VMSME_L3PHIC20n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(3),
        VMSME_L3PHIC20n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(3),
        VMSME_L3PHIC20n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(3),
        VMSME_L3PHIC20n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(3),
        VMSME_L3PHIC20n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(3),
        VMSME_L3PHIC20n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(3),
        VMSME_L3PHIC20n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(3),
        VMSME_L3PHIC20n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(3),
        VMSME_L3PHIC20n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(3),
        VMSME_L3PHIC20n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(3),
        VMSME_L3PHIC20n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(3),
        VMSME_L3PHIC20n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(3),
        VMSME_L3PHIC20n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(3),
        VMSME_L3PHIC20n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(3),
        VMSME_L3PHIC20n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(3),
        VMSME_L3PHIC20n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(3),
        VMSME_L3PHIC20n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(3),
        VMSME_L3PHIC20n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(3),
        VMSME_L3PHIC20n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(3),
        VMSME_L3PHIC20n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(3),
        VMSME_L3PHIC20n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(3),
        VMSME_L3PHIC20n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(3),
        VMSME_L3PHIC20n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(3),
        VMSME_L3PHIC20n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(3),
        VMSME_L3PHIC20n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(3),
        VMSME_L3PHIC20n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(3),
        VMSME_L3PHIC20n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(3),
        VMSME_L3PHIC20n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(3),
        VMSME_L3PHIC20n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(3),
        VMSME_L3PHIC20n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(3),
        VMSME_L3PHIC20n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(3),
        VMSME_L3PHIC20n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(3),
        VMSME_L3PHIC20n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(3),
        VMSME_L3PHIC20n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(3),
        VMSME_L3PHIC20n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(3),
        VMSME_L3PHIC20n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(3),
        VMSME_L3PHIC20n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(3),
        VMSME_L3PHIC20n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(3),
        VMSME_L3PHIC20n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(3),
        VMSME_L3PHIC20n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(3),
        VMSME_L3PHIC20n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(3),
        VMSME_L3PHIC20n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(3),
        VMSME_L3PHIC20n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(3),
        VMSME_L3PHIC20n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(3),
        VMSME_L3PHIC20n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(3),
        VMSME_L3PHIC20n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(3),
        VMSME_L3PHIC20n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(3),
        VMSME_L3PHIC20n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(3),
        VMSME_L3PHIC20n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(3),
        VMSME_L3PHIC20n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(3),
        VMSME_L3PHIC20n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(3),
        VMSME_L3PHIC20n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(3),
        VMSME_L3PHIC20n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(3),
        VMSME_L3PHIC20n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(3),
        VMSME_L3PHIC20n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(3),
        VMSME_L3PHIC20n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(3),
        VMSME_L3PHIC20n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(3),
        VMSME_L3PHIC20n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(3),
        VMSME_L3PHIC20n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(3),
        VMSME_L3PHIC20n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(3),
        VMSME_L3PHIC20n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(3),
        VMSME_L3PHIC20n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(3),
        VMSME_L3PHIC20n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(3),
        VMSME_L3PHIC20n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(3),
        VMSME_L3PHIC20n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(3),
        VMSME_L3PHIC20n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(3),
        VMSME_L3PHIC20n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(3),
        VMSME_L3PHIC20n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(3),
        VMSME_L3PHIC20n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(3),
        VMSME_L3PHIC20n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(3),
        VMSME_L3PHIC20n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(3),
        VMSME_L3PHIC20n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(3),
        VMSME_L3PHIC20n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(3),
        VMSME_L3PHIC21n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(4),
        VMSME_L3PHIC21n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(4),
        VMSME_L3PHIC21n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(4),
        VMSME_L3PHIC21n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(4),
        VMSME_L3PHIC21n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(4),
        VMSME_L3PHIC21n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(4),
        VMSME_L3PHIC21n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(4),
        VMSME_L3PHIC21n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(4),
        VMSME_L3PHIC21n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(4),
        VMSME_L3PHIC21n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(4),
        VMSME_L3PHIC21n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(4),
        VMSME_L3PHIC21n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(4),
        VMSME_L3PHIC21n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(4),
        VMSME_L3PHIC21n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(4),
        VMSME_L3PHIC21n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(4),
        VMSME_L3PHIC21n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(4),
        VMSME_L3PHIC21n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(4),
        VMSME_L3PHIC21n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(4),
        VMSME_L3PHIC21n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(4),
        VMSME_L3PHIC21n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(4),
        VMSME_L3PHIC21n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(4),
        VMSME_L3PHIC21n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(4),
        VMSME_L3PHIC21n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(4),
        VMSME_L3PHIC21n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(4),
        VMSME_L3PHIC21n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(4),
        VMSME_L3PHIC21n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(4),
        VMSME_L3PHIC21n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(4),
        VMSME_L3PHIC21n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(4),
        VMSME_L3PHIC21n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(4),
        VMSME_L3PHIC21n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(4),
        VMSME_L3PHIC21n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(4),
        VMSME_L3PHIC21n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(4),
        VMSME_L3PHIC21n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(4),
        VMSME_L3PHIC21n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(4),
        VMSME_L3PHIC21n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(4),
        VMSME_L3PHIC21n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(4),
        VMSME_L3PHIC21n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(4),
        VMSME_L3PHIC21n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(4),
        VMSME_L3PHIC21n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(4),
        VMSME_L3PHIC21n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(4),
        VMSME_L3PHIC21n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(4),
        VMSME_L3PHIC21n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(4),
        VMSME_L3PHIC21n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(4),
        VMSME_L3PHIC21n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(4),
        VMSME_L3PHIC21n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(4),
        VMSME_L3PHIC21n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(4),
        VMSME_L3PHIC21n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(4),
        VMSME_L3PHIC21n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(4),
        VMSME_L3PHIC21n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(4),
        VMSME_L3PHIC21n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(4),
        VMSME_L3PHIC21n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(4),
        VMSME_L3PHIC21n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(4),
        VMSME_L3PHIC21n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(4),
        VMSME_L3PHIC21n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(4),
        VMSME_L3PHIC21n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(4),
        VMSME_L3PHIC21n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(4),
        VMSME_L3PHIC21n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(4),
        VMSME_L3PHIC21n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(4),
        VMSME_L3PHIC21n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(4),
        VMSME_L3PHIC21n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(4),
        VMSME_L3PHIC21n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(4),
        VMSME_L3PHIC21n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(4),
        VMSME_L3PHIC21n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(4),
        VMSME_L3PHIC21n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(4),
        VMSME_L3PHIC21n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(4),
        VMSME_L3PHIC21n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(4),
        VMSME_L3PHIC21n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(4),
        VMSME_L3PHIC21n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(4),
        VMSME_L3PHIC21n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(4),
        VMSME_L3PHIC21n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(4),
        VMSME_L3PHIC21n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(4),
        VMSME_L3PHIC21n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(4),
        VMSME_L3PHIC21n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(4),
        VMSME_L3PHIC21n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(4),
        VMSME_L3PHIC21n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(4),
        VMSME_L3PHIC21n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(4),
        VMSME_L3PHIC21n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(4),
        VMSME_L3PHIC21n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(4),
        VMSME_L3PHIC21n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(4),
        VMSME_L3PHIC21n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(4),
        VMSME_L3PHIC21n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(4),
        VMSME_L3PHIC21n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(4),
        VMSME_L3PHIC21n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(4),
        VMSME_L3PHIC21n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(4),
        VMSME_L3PHIC21n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(4),
        VMSME_L3PHIC21n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(4),
        VMSME_L3PHIC21n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(4),
        VMSME_L3PHIC21n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(4),
        VMSME_L3PHIC21n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(4),
        VMSME_L3PHIC21n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(4),
        VMSME_L3PHIC21n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(4),
        VMSME_L3PHIC21n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(4),
        VMSME_L3PHIC21n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(4),
        VMSME_L3PHIC21n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(4),
        VMSME_L3PHIC21n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(4),
        VMSME_L3PHIC21n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(4),
        VMSME_L3PHIC21n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(4),
        VMSME_L3PHIC21n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(4),
        VMSME_L3PHIC21n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(4),
        VMSME_L3PHIC21n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(4),
        VMSME_L3PHIC21n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(4),
        VMSME_L3PHIC21n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(4),
        VMSME_L3PHIC21n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(4),
        VMSME_L3PHIC21n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(4),
        VMSME_L3PHIC21n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(4),
        VMSME_L3PHIC21n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(4),
        VMSME_L3PHIC21n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(4),
        VMSME_L3PHIC21n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(4),
        VMSME_L3PHIC21n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(4),
        VMSME_L3PHIC21n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(4),
        VMSME_L3PHIC21n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(4),
        VMSME_L3PHIC21n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(4),
        VMSME_L3PHIC21n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(4),
        VMSME_L3PHIC21n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(4),
        VMSME_L3PHIC21n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(4),
        VMSME_L3PHIC21n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(4),
        VMSME_L3PHIC21n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(4),
        VMSME_L3PHIC21n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(4),
        VMSME_L3PHIC21n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(4),
        VMSME_L3PHIC21n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(4),
        VMSME_L3PHIC21n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(4),
        VMSME_L3PHIC21n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(4),
        VMSME_L3PHIC21n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(4),
        VMSME_L3PHIC21n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(4),
        VMSME_L3PHIC21n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(4),
        VMSME_L3PHIC21n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(4),
        VMSME_L3PHIC21n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(4),
        VMSME_L3PHIC21n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(4),
        VMSME_L3PHIC21n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(4),
        VMSME_L3PHIC21n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(4),
        VMSME_L3PHIC21n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(4),
        VMSME_L3PHIC22n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(5),
        VMSME_L3PHIC22n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(5),
        VMSME_L3PHIC22n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(5),
        VMSME_L3PHIC22n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(5),
        VMSME_L3PHIC22n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(5),
        VMSME_L3PHIC22n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(5),
        VMSME_L3PHIC22n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(5),
        VMSME_L3PHIC22n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(5),
        VMSME_L3PHIC22n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(5),
        VMSME_L3PHIC22n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(5),
        VMSME_L3PHIC22n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(5),
        VMSME_L3PHIC22n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(5),
        VMSME_L3PHIC22n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(5),
        VMSME_L3PHIC22n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(5),
        VMSME_L3PHIC22n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(5),
        VMSME_L3PHIC22n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(5),
        VMSME_L3PHIC22n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(5),
        VMSME_L3PHIC22n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(5),
        VMSME_L3PHIC22n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(5),
        VMSME_L3PHIC22n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(5),
        VMSME_L3PHIC22n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(5),
        VMSME_L3PHIC22n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(5),
        VMSME_L3PHIC22n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(5),
        VMSME_L3PHIC22n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(5),
        VMSME_L3PHIC22n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(5),
        VMSME_L3PHIC22n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(5),
        VMSME_L3PHIC22n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(5),
        VMSME_L3PHIC22n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(5),
        VMSME_L3PHIC22n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(5),
        VMSME_L3PHIC22n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(5),
        VMSME_L3PHIC22n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(5),
        VMSME_L3PHIC22n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(5),
        VMSME_L3PHIC22n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(5),
        VMSME_L3PHIC22n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(5),
        VMSME_L3PHIC22n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(5),
        VMSME_L3PHIC22n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(5),
        VMSME_L3PHIC22n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(5),
        VMSME_L3PHIC22n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(5),
        VMSME_L3PHIC22n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(5),
        VMSME_L3PHIC22n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(5),
        VMSME_L3PHIC22n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(5),
        VMSME_L3PHIC22n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(5),
        VMSME_L3PHIC22n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(5),
        VMSME_L3PHIC22n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(5),
        VMSME_L3PHIC22n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(5),
        VMSME_L3PHIC22n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(5),
        VMSME_L3PHIC22n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(5),
        VMSME_L3PHIC22n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(5),
        VMSME_L3PHIC22n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(5),
        VMSME_L3PHIC22n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(5),
        VMSME_L3PHIC22n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(5),
        VMSME_L3PHIC22n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(5),
        VMSME_L3PHIC22n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(5),
        VMSME_L3PHIC22n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(5),
        VMSME_L3PHIC22n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(5),
        VMSME_L3PHIC22n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(5),
        VMSME_L3PHIC22n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(5),
        VMSME_L3PHIC22n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(5),
        VMSME_L3PHIC22n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(5),
        VMSME_L3PHIC22n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(5),
        VMSME_L3PHIC22n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(5),
        VMSME_L3PHIC22n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(5),
        VMSME_L3PHIC22n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(5),
        VMSME_L3PHIC22n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(5),
        VMSME_L3PHIC22n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(5),
        VMSME_L3PHIC22n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(5),
        VMSME_L3PHIC22n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(5),
        VMSME_L3PHIC22n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(5),
        VMSME_L3PHIC22n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(5),
        VMSME_L3PHIC22n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(5),
        VMSME_L3PHIC22n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(5),
        VMSME_L3PHIC22n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(5),
        VMSME_L3PHIC22n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(5),
        VMSME_L3PHIC22n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(5),
        VMSME_L3PHIC22n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(5),
        VMSME_L3PHIC22n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(5),
        VMSME_L3PHIC22n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(5),
        VMSME_L3PHIC22n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(5),
        VMSME_L3PHIC22n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(5),
        VMSME_L3PHIC22n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(5),
        VMSME_L3PHIC22n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(5),
        VMSME_L3PHIC22n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(5),
        VMSME_L3PHIC22n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(5),
        VMSME_L3PHIC22n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(5),
        VMSME_L3PHIC22n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(5),
        VMSME_L3PHIC22n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(5),
        VMSME_L3PHIC22n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(5),
        VMSME_L3PHIC22n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(5),
        VMSME_L3PHIC22n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(5),
        VMSME_L3PHIC22n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(5),
        VMSME_L3PHIC22n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(5),
        VMSME_L3PHIC22n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(5),
        VMSME_L3PHIC22n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(5),
        VMSME_L3PHIC22n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(5),
        VMSME_L3PHIC22n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(5),
        VMSME_L3PHIC22n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(5),
        VMSME_L3PHIC22n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(5),
        VMSME_L3PHIC22n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(5),
        VMSME_L3PHIC22n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(5),
        VMSME_L3PHIC22n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(5),
        VMSME_L3PHIC22n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(5),
        VMSME_L3PHIC22n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(5),
        VMSME_L3PHIC22n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(5),
        VMSME_L3PHIC22n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(5),
        VMSME_L3PHIC22n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(5),
        VMSME_L3PHIC22n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(5),
        VMSME_L3PHIC22n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(5),
        VMSME_L3PHIC22n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(5),
        VMSME_L3PHIC22n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(5),
        VMSME_L3PHIC22n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(5),
        VMSME_L3PHIC22n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(5),
        VMSME_L3PHIC22n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(5),
        VMSME_L3PHIC22n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(5),
        VMSME_L3PHIC22n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(5),
        VMSME_L3PHIC22n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(5),
        VMSME_L3PHIC22n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(5),
        VMSME_L3PHIC22n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(5),
        VMSME_L3PHIC22n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(5),
        VMSME_L3PHIC22n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(5),
        VMSME_L3PHIC22n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(5),
        VMSME_L3PHIC22n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(5),
        VMSME_L3PHIC22n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(5),
        VMSME_L3PHIC22n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(5),
        VMSME_L3PHIC22n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(5),
        VMSME_L3PHIC22n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(5),
        VMSME_L3PHIC22n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(5),
        VMSME_L3PHIC22n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(5),
        VMSME_L3PHIC22n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(5),
        VMSME_L3PHIC22n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(5),
        VMSME_L3PHIC22n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(5),
        VMSME_L3PHIC22n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(5),
        VMSME_L3PHIC23n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(6),
        VMSME_L3PHIC23n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(6),
        VMSME_L3PHIC23n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(6),
        VMSME_L3PHIC23n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(6),
        VMSME_L3PHIC23n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(6),
        VMSME_L3PHIC23n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(6),
        VMSME_L3PHIC23n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(6),
        VMSME_L3PHIC23n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(6),
        VMSME_L3PHIC23n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(6),
        VMSME_L3PHIC23n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(6),
        VMSME_L3PHIC23n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(6),
        VMSME_L3PHIC23n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(6),
        VMSME_L3PHIC23n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(6),
        VMSME_L3PHIC23n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(6),
        VMSME_L3PHIC23n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(6),
        VMSME_L3PHIC23n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(6),
        VMSME_L3PHIC23n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(6),
        VMSME_L3PHIC23n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(6),
        VMSME_L3PHIC23n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(6),
        VMSME_L3PHIC23n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(6),
        VMSME_L3PHIC23n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(6),
        VMSME_L3PHIC23n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(6),
        VMSME_L3PHIC23n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(6),
        VMSME_L3PHIC23n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(6),
        VMSME_L3PHIC23n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(6),
        VMSME_L3PHIC23n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(6),
        VMSME_L3PHIC23n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(6),
        VMSME_L3PHIC23n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(6),
        VMSME_L3PHIC23n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(6),
        VMSME_L3PHIC23n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(6),
        VMSME_L3PHIC23n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(6),
        VMSME_L3PHIC23n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(6),
        VMSME_L3PHIC23n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(6),
        VMSME_L3PHIC23n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(6),
        VMSME_L3PHIC23n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(6),
        VMSME_L3PHIC23n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(6),
        VMSME_L3PHIC23n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(6),
        VMSME_L3PHIC23n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(6),
        VMSME_L3PHIC23n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(6),
        VMSME_L3PHIC23n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(6),
        VMSME_L3PHIC23n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(6),
        VMSME_L3PHIC23n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(6),
        VMSME_L3PHIC23n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(6),
        VMSME_L3PHIC23n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(6),
        VMSME_L3PHIC23n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(6),
        VMSME_L3PHIC23n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(6),
        VMSME_L3PHIC23n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(6),
        VMSME_L3PHIC23n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(6),
        VMSME_L3PHIC23n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(6),
        VMSME_L3PHIC23n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(6),
        VMSME_L3PHIC23n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(6),
        VMSME_L3PHIC23n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(6),
        VMSME_L3PHIC23n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(6),
        VMSME_L3PHIC23n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(6),
        VMSME_L3PHIC23n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(6),
        VMSME_L3PHIC23n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(6),
        VMSME_L3PHIC23n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(6),
        VMSME_L3PHIC23n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(6),
        VMSME_L3PHIC23n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(6),
        VMSME_L3PHIC23n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(6),
        VMSME_L3PHIC23n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(6),
        VMSME_L3PHIC23n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(6),
        VMSME_L3PHIC23n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(6),
        VMSME_L3PHIC23n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(6),
        VMSME_L3PHIC23n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(6),
        VMSME_L3PHIC23n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(6),
        VMSME_L3PHIC23n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(6),
        VMSME_L3PHIC23n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(6),
        VMSME_L3PHIC23n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(6),
        VMSME_L3PHIC23n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(6),
        VMSME_L3PHIC23n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(6),
        VMSME_L3PHIC23n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(6),
        VMSME_L3PHIC23n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(6),
        VMSME_L3PHIC23n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(6),
        VMSME_L3PHIC23n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(6),
        VMSME_L3PHIC23n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(6),
        VMSME_L3PHIC23n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(6),
        VMSME_L3PHIC23n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(6),
        VMSME_L3PHIC23n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(6),
        VMSME_L3PHIC23n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(6),
        VMSME_L3PHIC23n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(6),
        VMSME_L3PHIC23n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(6),
        VMSME_L3PHIC23n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(6),
        VMSME_L3PHIC23n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(6),
        VMSME_L3PHIC23n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(6),
        VMSME_L3PHIC23n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(6),
        VMSME_L3PHIC23n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(6),
        VMSME_L3PHIC23n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(6),
        VMSME_L3PHIC23n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(6),
        VMSME_L3PHIC23n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(6),
        VMSME_L3PHIC23n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(6),
        VMSME_L3PHIC23n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(6),
        VMSME_L3PHIC23n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(6),
        VMSME_L3PHIC23n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(6),
        VMSME_L3PHIC23n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(6),
        VMSME_L3PHIC23n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(6),
        VMSME_L3PHIC23n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(6),
        VMSME_L3PHIC23n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(6),
        VMSME_L3PHIC23n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(6),
        VMSME_L3PHIC23n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(6),
        VMSME_L3PHIC23n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(6),
        VMSME_L3PHIC23n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(6),
        VMSME_L3PHIC23n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(6),
        VMSME_L3PHIC23n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(6),
        VMSME_L3PHIC23n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(6),
        VMSME_L3PHIC23n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(6),
        VMSME_L3PHIC23n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(6),
        VMSME_L3PHIC23n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(6),
        VMSME_L3PHIC23n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(6),
        VMSME_L3PHIC23n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(6),
        VMSME_L3PHIC23n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(6),
        VMSME_L3PHIC23n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(6),
        VMSME_L3PHIC23n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(6),
        VMSME_L3PHIC23n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(6),
        VMSME_L3PHIC23n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(6),
        VMSME_L3PHIC23n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(6),
        VMSME_L3PHIC23n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(6),
        VMSME_L3PHIC23n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(6),
        VMSME_L3PHIC23n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(6),
        VMSME_L3PHIC23n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(6),
        VMSME_L3PHIC23n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(6),
        VMSME_L3PHIC23n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(6),
        VMSME_L3PHIC23n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(6),
        VMSME_L3PHIC23n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(6),
        VMSME_L3PHIC23n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(6),
        VMSME_L3PHIC23n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(6),
        VMSME_L3PHIC23n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(6),
        VMSME_L3PHIC23n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(6),
        VMSME_L3PHIC23n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(6),
        VMSME_L3PHIC23n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(6),
        VMSME_L3PHIC23n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(6),
        VMSME_L3PHIC24n1_dataarray_data_V_wea       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_wea(7),
        VMSME_L3PHIC24n1_dataarray_data_V_writeaddr => VMSME_L3PHIC17to24n1_dataarray_data_V_writeaddr(7),
        VMSME_L3PHIC24n1_dataarray_data_V_din       =>       VMSME_L3PHIC17to24n1_dataarray_data_V_din(7),
        VMSME_L3PHIC24n1_nentries_0_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(0)(7),
        VMSME_L3PHIC24n1_nentries_0_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(0)(7),
        VMSME_L3PHIC24n1_nentries_0_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(1)(7),
        VMSME_L3PHIC24n1_nentries_0_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(1)(7),
        VMSME_L3PHIC24n1_nentries_0_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(2)(7),
        VMSME_L3PHIC24n1_nentries_0_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(2)(7),
        VMSME_L3PHIC24n1_nentries_0_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(3)(7),
        VMSME_L3PHIC24n1_nentries_0_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(3)(7),
        VMSME_L3PHIC24n1_nentries_0_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(4)(7),
        VMSME_L3PHIC24n1_nentries_0_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(4)(7),
        VMSME_L3PHIC24n1_nentries_0_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(5)(7),
        VMSME_L3PHIC24n1_nentries_0_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(5)(7),
        VMSME_L3PHIC24n1_nentries_0_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(6)(7),
        VMSME_L3PHIC24n1_nentries_0_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(6)(7),
        VMSME_L3PHIC24n1_nentries_0_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(0)(7)(7),
        VMSME_L3PHIC24n1_nentries_0_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(0)(7)(7),
        VMSME_L3PHIC24n1_nentries_1_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(0)(7),
        VMSME_L3PHIC24n1_nentries_1_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(0)(7),
        VMSME_L3PHIC24n1_nentries_1_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(1)(7),
        VMSME_L3PHIC24n1_nentries_1_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(1)(7),
        VMSME_L3PHIC24n1_nentries_1_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(2)(7),
        VMSME_L3PHIC24n1_nentries_1_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(2)(7),
        VMSME_L3PHIC24n1_nentries_1_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(3)(7),
        VMSME_L3PHIC24n1_nentries_1_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(3)(7),
        VMSME_L3PHIC24n1_nentries_1_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(4)(7),
        VMSME_L3PHIC24n1_nentries_1_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(4)(7),
        VMSME_L3PHIC24n1_nentries_1_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(5)(7),
        VMSME_L3PHIC24n1_nentries_1_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(5)(7),
        VMSME_L3PHIC24n1_nentries_1_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(6)(7),
        VMSME_L3PHIC24n1_nentries_1_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(6)(7),
        VMSME_L3PHIC24n1_nentries_1_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(1)(7)(7),
        VMSME_L3PHIC24n1_nentries_1_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(1)(7)(7),
        VMSME_L3PHIC24n1_nentries_2_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(0)(7),
        VMSME_L3PHIC24n1_nentries_2_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(0)(7),
        VMSME_L3PHIC24n1_nentries_2_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(1)(7),
        VMSME_L3PHIC24n1_nentries_2_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(1)(7),
        VMSME_L3PHIC24n1_nentries_2_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(2)(7),
        VMSME_L3PHIC24n1_nentries_2_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(2)(7),
        VMSME_L3PHIC24n1_nentries_2_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(3)(7),
        VMSME_L3PHIC24n1_nentries_2_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(3)(7),
        VMSME_L3PHIC24n1_nentries_2_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(4)(7),
        VMSME_L3PHIC24n1_nentries_2_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(4)(7),
        VMSME_L3PHIC24n1_nentries_2_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(5)(7),
        VMSME_L3PHIC24n1_nentries_2_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(5)(7),
        VMSME_L3PHIC24n1_nentries_2_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(6)(7),
        VMSME_L3PHIC24n1_nentries_2_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(6)(7),
        VMSME_L3PHIC24n1_nentries_2_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(2)(7)(7),
        VMSME_L3PHIC24n1_nentries_2_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(2)(7)(7),
        VMSME_L3PHIC24n1_nentries_3_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(0)(7),
        VMSME_L3PHIC24n1_nentries_3_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(0)(7),
        VMSME_L3PHIC24n1_nentries_3_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(1)(7),
        VMSME_L3PHIC24n1_nentries_3_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(1)(7),
        VMSME_L3PHIC24n1_nentries_3_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(2)(7),
        VMSME_L3PHIC24n1_nentries_3_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(2)(7),
        VMSME_L3PHIC24n1_nentries_3_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(3)(7),
        VMSME_L3PHIC24n1_nentries_3_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(3)(7),
        VMSME_L3PHIC24n1_nentries_3_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(4)(7),
        VMSME_L3PHIC24n1_nentries_3_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(4)(7),
        VMSME_L3PHIC24n1_nentries_3_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(5)(7),
        VMSME_L3PHIC24n1_nentries_3_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(5)(7),
        VMSME_L3PHIC24n1_nentries_3_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(6)(7),
        VMSME_L3PHIC24n1_nentries_3_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(6)(7),
        VMSME_L3PHIC24n1_nentries_3_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(3)(7)(7),
        VMSME_L3PHIC24n1_nentries_3_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(3)(7)(7),
        VMSME_L3PHIC24n1_nentries_4_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(0)(7),
        VMSME_L3PHIC24n1_nentries_4_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(0)(7),
        VMSME_L3PHIC24n1_nentries_4_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(1)(7),
        VMSME_L3PHIC24n1_nentries_4_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(1)(7),
        VMSME_L3PHIC24n1_nentries_4_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(2)(7),
        VMSME_L3PHIC24n1_nentries_4_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(2)(7),
        VMSME_L3PHIC24n1_nentries_4_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(3)(7),
        VMSME_L3PHIC24n1_nentries_4_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(3)(7),
        VMSME_L3PHIC24n1_nentries_4_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(4)(7),
        VMSME_L3PHIC24n1_nentries_4_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(4)(7),
        VMSME_L3PHIC24n1_nentries_4_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(5)(7),
        VMSME_L3PHIC24n1_nentries_4_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(5)(7),
        VMSME_L3PHIC24n1_nentries_4_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(6)(7),
        VMSME_L3PHIC24n1_nentries_4_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(6)(7),
        VMSME_L3PHIC24n1_nentries_4_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(4)(7)(7),
        VMSME_L3PHIC24n1_nentries_4_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(4)(7)(7),
        VMSME_L3PHIC24n1_nentries_5_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(0)(7),
        VMSME_L3PHIC24n1_nentries_5_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(0)(7),
        VMSME_L3PHIC24n1_nentries_5_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(1)(7),
        VMSME_L3PHIC24n1_nentries_5_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(1)(7),
        VMSME_L3PHIC24n1_nentries_5_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(2)(7),
        VMSME_L3PHIC24n1_nentries_5_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(2)(7),
        VMSME_L3PHIC24n1_nentries_5_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(3)(7),
        VMSME_L3PHIC24n1_nentries_5_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(3)(7),
        VMSME_L3PHIC24n1_nentries_5_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(4)(7),
        VMSME_L3PHIC24n1_nentries_5_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(4)(7),
        VMSME_L3PHIC24n1_nentries_5_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(5)(7),
        VMSME_L3PHIC24n1_nentries_5_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(5)(7),
        VMSME_L3PHIC24n1_nentries_5_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(6)(7),
        VMSME_L3PHIC24n1_nentries_5_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(6)(7),
        VMSME_L3PHIC24n1_nentries_5_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(5)(7)(7),
        VMSME_L3PHIC24n1_nentries_5_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(5)(7)(7),
        VMSME_L3PHIC24n1_nentries_6_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(0)(7),
        VMSME_L3PHIC24n1_nentries_6_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(0)(7),
        VMSME_L3PHIC24n1_nentries_6_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(1)(7),
        VMSME_L3PHIC24n1_nentries_6_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(1)(7),
        VMSME_L3PHIC24n1_nentries_6_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(2)(7),
        VMSME_L3PHIC24n1_nentries_6_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(2)(7),
        VMSME_L3PHIC24n1_nentries_6_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(3)(7),
        VMSME_L3PHIC24n1_nentries_6_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(3)(7),
        VMSME_L3PHIC24n1_nentries_6_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(4)(7),
        VMSME_L3PHIC24n1_nentries_6_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(4)(7),
        VMSME_L3PHIC24n1_nentries_6_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(5)(7),
        VMSME_L3PHIC24n1_nentries_6_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(5)(7),
        VMSME_L3PHIC24n1_nentries_6_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(6)(7),
        VMSME_L3PHIC24n1_nentries_6_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(6)(7),
        VMSME_L3PHIC24n1_nentries_6_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(6)(7)(7),
        VMSME_L3PHIC24n1_nentries_6_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(6)(7)(7),
        VMSME_L3PHIC24n1_nentries_7_V_0_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(0)(7),
        VMSME_L3PHIC24n1_nentries_7_V_0_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(0)(7),
        VMSME_L3PHIC24n1_nentries_7_V_1_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(1)(7),
        VMSME_L3PHIC24n1_nentries_7_V_1_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(1)(7),
        VMSME_L3PHIC24n1_nentries_7_V_2_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(2)(7),
        VMSME_L3PHIC24n1_nentries_7_V_2_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(2)(7),
        VMSME_L3PHIC24n1_nentries_7_V_3_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(3)(7),
        VMSME_L3PHIC24n1_nentries_7_V_3_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(3)(7),
        VMSME_L3PHIC24n1_nentries_7_V_4_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(4)(7),
        VMSME_L3PHIC24n1_nentries_7_V_4_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(4)(7),
        VMSME_L3PHIC24n1_nentries_7_V_5_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(5)(7),
        VMSME_L3PHIC24n1_nentries_7_V_5_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(5)(7),
        VMSME_L3PHIC24n1_nentries_7_V_6_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(6)(7),
        VMSME_L3PHIC24n1_nentries_7_V_6_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(6)(7),
        VMSME_L3PHIC24n1_nentries_7_V_7_we  =>  VMSME_L3PHIC17to24n1_nentries_V_we(7)(7)(7),
        VMSME_L3PHIC24n1_nentries_7_V_7_din => VMSME_L3PHIC17to24n1_nentries_V_din(7)(7)(7),
        AS_L3PHICn6_dataarray_data_V_wea       => AS_L3PHICn4_dataarray_data_V_wea,
        AS_L3PHICn6_dataarray_data_V_writeaddr => AS_L3PHICn4_dataarray_data_V_writeaddr,
        AS_L3PHICn6_dataarray_data_V_din       => AS_L3PHICn4_dataarray_data_V_din,
        AS_L3PHICn6_nentries_0_V_we  =>  AS_L3PHICn4_nentries_V_we(0),
        AS_L3PHICn6_nentries_0_V_din => AS_L3PHICn4_nentries_V_din(0),
        AS_L3PHICn6_nentries_1_V_we  =>  AS_L3PHICn4_nentries_V_we(1),
        AS_L3PHICn6_nentries_1_V_din => AS_L3PHICn4_nentries_V_din(1),
        AS_L3PHICn6_nentries_2_V_we  =>  AS_L3PHICn4_nentries_V_we(2),
        AS_L3PHICn6_nentries_2_V_din => AS_L3PHICn4_nentries_V_din(2),
        AS_L3PHICn6_nentries_3_V_we  =>  AS_L3PHICn4_nentries_V_we(3),
        AS_L3PHICn6_nentries_3_V_din => AS_L3PHICn4_nentries_V_din(3),
        AS_L3PHICn6_nentries_4_V_we  =>  AS_L3PHICn4_nentries_V_we(4),
        AS_L3PHICn6_nentries_4_V_din => AS_L3PHICn4_nentries_V_din(4),
        AS_L3PHICn6_nentries_5_V_we  =>  AS_L3PHICn4_nentries_V_we(5),
        AS_L3PHICn6_nentries_5_V_din => AS_L3PHICn4_nentries_V_din(5),
        AS_L3PHICn6_nentries_6_V_we  =>  AS_L3PHICn4_nentries_V_we(6),
        AS_L3PHICn6_nentries_6_V_din => AS_L3PHICn4_nentries_V_din(6),
        AS_L3PHICn6_nentries_7_V_we  =>  AS_L3PHICn4_nentries_V_we(7),
        AS_L3PHICn6_nentries_7_V_din => AS_L3PHICn4_nentries_V_din(7),
        FM_L1L2XX_L3PHIC_dataarray_data_V_enb      => FM_L1L2XX_L3PHIC_dataarray_data_V_enb,
        FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr => FM_L1L2XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L1L2XX_L3PHIC_dataarray_data_V_dout     => FM_L1L2XX_L3PHIC_dataarray_data_V_dout,
        FM_L1L2XX_L3PHIC_nentries_0_V_dout         => FM_L1L2XX_L3PHIC_nentries_V_dout(0),
        FM_L1L2XX_L3PHIC_nentries_1_V_dout         => FM_L1L2XX_L3PHIC_nentries_V_dout(1),
        FM_L5L6XX_L3PHIC_dataarray_data_V_enb      => FM_L5L6XX_L3PHIC_dataarray_data_V_enb,
        FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr => FM_L5L6XX_L3PHIC_dataarray_data_V_readaddr,
        FM_L5L6XX_L3PHIC_dataarray_data_V_dout     => FM_L5L6XX_L3PHIC_dataarray_data_V_dout,
        FM_L5L6XX_L3PHIC_nentries_0_V_dout         => FM_L5L6XX_L3PHIC_nentries_V_dout(0),
        FM_L5L6XX_L3PHIC_nentries_1_V_dout         => FM_L5L6XX_L3PHIC_nentries_V_dout(1)  );
  end generate;


end behavior;
