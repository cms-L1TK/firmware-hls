-------------------------------------------------------------------------------
-- Title      : tf wrapper
-- Project    : 
-------------------------------------------------------------------------------
-- File       : tf_wrapper.vhd
-- Author     : Michael Oshiro  <mco62@cornell.edu>
-- Company    : Cornell University
-- Created    : 2024-01-19
-- Last update: 2024-01-19
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Simple module to pack/unpack SectorProcessor inputs into vectors
-------------------------------------------------------------------------------
-- Copyright (c) 2024 Cornell University
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2022-01-19  1.0      oshiro  Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

use work.memUtil_pkg.all;
use work.memUtil_aux_pkg_f2.all;

entity tf2_wrapper is
  port (
    clk                       : in  std_logic;
    reset                     : in  std_logic;
    start_first_write         : in  std_logic;
    PC_start                  : in  std_logic;
    PC_bx_in                  : in  std_logic_vector(2 downto 0);
    FT_bx_out_0               : out std_logic_vector(2 downto 0); 
    FT_bx_out_vld             : out std_logic;
    FT_done                   : out std_logic;
    FT_last_track             : out std_logic;
    FT_last_track_vld         : out std_logic;
    AS_36_wea                 : in t_arr_AS_36_1b;
    AS_36_writeaddr           : in t_arr_AS_36_ADDR;
    AS_36_din                 : in t_arr_AS_36_DATA;
    MPAR_73_wea               : in t_arr_MTPAR_73_1b;
    MPAR_73_writeaddr         : in t_arr_MTPAR_73_ADDR;
    MPAR_73_din               : in t_arr_MTPAR_73_DATA;
    TW_104_stream_AV_din      : out t_arr_TW_104_DATA;
    TW_104_stream_A_full_neg  : in t_arr_TW_104_1b;
    TW_104_stream_A_write     : out t_arr_TW_104_1b;
    DW_49_stream_AV_din       : out t_arr_DW_49_DATA;
    DW_49_stream_A_full_neg   : in t_arr_DW_49_1b;
    DW_49_stream_A_write      : out t_arr_DW_49_1b;
    BW_46_stream_AV_din       : out t_arr_BW_46_DATA;
    BW_46_stream_A_full_neg   : in t_arr_BW_46_1b;
    BW_46_stream_A_write      : out t_arr_BW_46_1b
    );
end entity tf2_wrapper;

architecture rtl of tf2_wrapper is

begin  -- architecture rtl

  SectorProcessor_1 : entity work.SectorProcessor
    port map (
      clk                     => clk,
      reset                   => reset,
      start_first_write       => start_first_write,
      PC_start                => PC_start,
      PC_bx_in                => PC_bx_in,
      FT_bx_out_0             => FT_bx_out_0,
      FT_bx_out_vld           => FT_bx_out_vld,
      FT_done                 => FT_done,
      FT_L1L2_last_track      => FT_last_track,
      FT_L1L2_last_track_vld  => FT_last_track_vld,
      FT_L2L3_last_track      => open,
      FT_L2L3_last_track_vld  => open,
      FT_L3L4_last_track      => open,
      FT_L3L4_last_track_vld  => open,
      FT_L5L6_last_track      => open,
      FT_L5L6_last_track_vld  => open,
      FT_D1D2_last_track      => open,
      FT_D1D2_last_track_vld  => open,
      FT_D3D4_last_track      => open,
      FT_D3D4_last_track_vld  => open,
      FT_L1D1_last_track      => open,
      FT_L1D1_last_track_vld  => open,
      FT_L2D1_last_track      => open,
      FT_L2D1_last_track_vld  => open,
      AS_L1PHIAin_wea       => AS_36_wea(L1PHIAn1),
      AS_L1PHIAin_writeaddr => AS_36_writeaddr(L1PHIAn1),
      AS_L1PHIAin_din       => AS_36_din(L1PHIAn1),
      AS_L1PHIBin_wea       => AS_36_wea(L1PHIBn1),
      AS_L1PHIBin_writeaddr => AS_36_writeaddr(L1PHIBn1),
      AS_L1PHIBin_din       => AS_36_din(L1PHIBn1),
      AS_L1PHICin_wea       => AS_36_wea(L1PHICn1),
      AS_L1PHICin_writeaddr => AS_36_writeaddr(L1PHICn1),
      AS_L1PHICin_din       => AS_36_din(L1PHICn1),
      AS_L1PHIDin_wea       => AS_36_wea(L1PHIDn1),
      AS_L1PHIDin_writeaddr => AS_36_writeaddr(L1PHIDn1),
      AS_L1PHIDin_din       => AS_36_din(L1PHIDn1),
      AS_L1PHIEin_wea       => AS_36_wea(L1PHIEn1),
      AS_L1PHIEin_writeaddr => AS_36_writeaddr(L1PHIEn1),
      AS_L1PHIEin_din       => AS_36_din(L1PHIEn1),
      AS_L1PHIFin_wea       => AS_36_wea(L1PHIFn1),
      AS_L1PHIFin_writeaddr => AS_36_writeaddr(L1PHIFn1),
      AS_L1PHIFin_din       => AS_36_din(L1PHIFn1),
      AS_L1PHIGin_wea       => AS_36_wea(L1PHIGn1),
      AS_L1PHIGin_writeaddr => AS_36_writeaddr(L1PHIGn1),
      AS_L1PHIGin_din       => AS_36_din(L1PHIGn1),
      AS_L1PHIHin_wea       => AS_36_wea(L1PHIHn1),
      AS_L1PHIHin_writeaddr => AS_36_writeaddr(L1PHIHn1),
      AS_L1PHIHin_din       => AS_36_din(L1PHIHn1),
      AS_L2PHIAin_wea       => AS_36_wea(L2PHIAn1),
      AS_L2PHIAin_writeaddr => AS_36_writeaddr(L2PHIAn1),
      AS_L2PHIAin_din       => AS_36_din(L2PHIAn1),
      AS_L2PHIBin_wea       => AS_36_wea(L2PHIBn1),
      AS_L2PHIBin_writeaddr => AS_36_writeaddr(L2PHIBn1),
      AS_L2PHIBin_din       => AS_36_din(L2PHIBn1),
      AS_L2PHICin_wea       => AS_36_wea(L2PHICn1),
      AS_L2PHICin_writeaddr => AS_36_writeaddr(L2PHICn1),
      AS_L2PHICin_din       => AS_36_din(L2PHICn1),
      AS_L2PHIDin_wea       => AS_36_wea(L2PHIDn1),
      AS_L2PHIDin_writeaddr => AS_36_writeaddr(L2PHIDn1),
      AS_L2PHIDin_din       => AS_36_din(L2PHIDn1),
      AS_L3PHIAin_wea       => AS_36_wea(L3PHIAn1),
      AS_L3PHIAin_writeaddr => AS_36_writeaddr(L3PHIAn1),
      AS_L3PHIAin_din       => AS_36_din(L3PHIAn1),
      AS_L3PHIBin_wea       => AS_36_wea(L3PHIBn1),
      AS_L3PHIBin_writeaddr => AS_36_writeaddr(L3PHIBn1),
      AS_L3PHIBin_din       => AS_36_din(L3PHIBn1),
      AS_L3PHICin_wea       => AS_36_wea(L3PHICn1),
      AS_L3PHICin_writeaddr => AS_36_writeaddr(L3PHICn1),
      AS_L3PHICin_din       => AS_36_din(L3PHICn1),
      AS_L3PHIDin_wea       => AS_36_wea(L3PHIDn1),
      AS_L3PHIDin_writeaddr => AS_36_writeaddr(L3PHIDn1),
      AS_L3PHIDin_din       => AS_36_din(L3PHIDn1),
      AS_L4PHIAin_wea       => AS_36_wea(L4PHIAn1),
      AS_L4PHIAin_writeaddr => AS_36_writeaddr(L4PHIAn1),
      AS_L4PHIAin_din       => AS_36_din(L4PHIAn1),
      AS_L4PHIBin_wea       => AS_36_wea(L4PHIBn1),
      AS_L4PHIBin_writeaddr => AS_36_writeaddr(L4PHIBn1),
      AS_L4PHIBin_din       => AS_36_din(L4PHIBn1),
      AS_L4PHICin_wea       => AS_36_wea(L4PHICn1),
      AS_L4PHICin_writeaddr => AS_36_writeaddr(L4PHICn1),
      AS_L4PHICin_din       => AS_36_din(L4PHICn1),
      AS_L4PHIDin_wea       => AS_36_wea(L4PHIDn1),
      AS_L4PHIDin_writeaddr => AS_36_writeaddr(L4PHIDn1),
      AS_L4PHIDin_din       => AS_36_din(L4PHIDn1),
      AS_L5PHIAin_wea       => AS_36_wea(L5PHIAn1),
      AS_L5PHIAin_writeaddr => AS_36_writeaddr(L5PHIAn1),
      AS_L5PHIAin_din       => AS_36_din(L5PHIAn1),
      AS_L5PHIBin_wea       => AS_36_wea(L5PHIBn1),
      AS_L5PHIBin_writeaddr => AS_36_writeaddr(L5PHIBn1),
      AS_L5PHIBin_din       => AS_36_din(L5PHIBn1),
      AS_L5PHICin_wea       => AS_36_wea(L5PHICn1),
      AS_L5PHICin_writeaddr => AS_36_writeaddr(L5PHICn1),
      AS_L5PHICin_din       => AS_36_din(L5PHICn1),
      AS_L5PHIDin_wea       => AS_36_wea(L5PHIDn1),
      AS_L5PHIDin_writeaddr => AS_36_writeaddr(L5PHIDn1),
      AS_L5PHIDin_din       => AS_36_din(L5PHIDn1),
      AS_L6PHIAin_wea       => AS_36_wea(L6PHIAn1),
      AS_L6PHIAin_writeaddr => AS_36_writeaddr(L6PHIAn1),
      AS_L6PHIAin_din       => AS_36_din(L6PHIAn1),
      AS_L6PHIBin_wea       => AS_36_wea(L6PHIBn1),
      AS_L6PHIBin_writeaddr => AS_36_writeaddr(L6PHIBn1),
      AS_L6PHIBin_din       => AS_36_din(L6PHIBn1),
      AS_L6PHICin_wea       => AS_36_wea(L6PHICn1),
      AS_L6PHICin_writeaddr => AS_36_writeaddr(L6PHICn1),
      AS_L6PHICin_din       => AS_36_din(L6PHICn1),
      AS_L6PHIDin_wea       => AS_36_wea(L6PHIDn1),
      AS_L6PHIDin_writeaddr => AS_36_writeaddr(L6PHIDn1),
      AS_L6PHIDin_din       => AS_36_din(L6PHIDn1),
      AS_D1PHIAin_wea       => AS_36_wea(D1PHIAn1),
      AS_D1PHIAin_writeaddr => AS_36_writeaddr(D1PHIAn1),
      AS_D1PHIAin_din       => AS_36_din(D1PHIAn1),
      AS_D1PHIBin_wea       => AS_36_wea(D1PHIBn1),
      AS_D1PHIBin_writeaddr => AS_36_writeaddr(D1PHIBn1),
      AS_D1PHIBin_din       => AS_36_din(D1PHIBn1),
      AS_D1PHICin_wea       => AS_36_wea(D1PHICn1),
      AS_D1PHICin_writeaddr => AS_36_writeaddr(D1PHICn1),
      AS_D1PHICin_din       => AS_36_din(D1PHICn1),
      AS_D1PHIDin_wea       => AS_36_wea(D1PHIDn1),
      AS_D1PHIDin_writeaddr => AS_36_writeaddr(D1PHIDn1),
      AS_D1PHIDin_din       => AS_36_din(D1PHIDn1),
      AS_D2PHIAin_wea       => AS_36_wea(D2PHIAn1),
      AS_D2PHIAin_writeaddr => AS_36_writeaddr(D2PHIAn1),
      AS_D2PHIAin_din       => AS_36_din(D2PHIAn1),
      AS_D2PHIBin_wea       => AS_36_wea(D2PHIBn1),
      AS_D2PHIBin_writeaddr => AS_36_writeaddr(D2PHIBn1),
      AS_D2PHIBin_din       => AS_36_din(D2PHIBn1),
      AS_D2PHICin_wea       => AS_36_wea(D2PHICn1),
      AS_D2PHICin_writeaddr => AS_36_writeaddr(D2PHICn1),
      AS_D2PHICin_din       => AS_36_din(D2PHICn1),
      AS_D2PHIDin_wea       => AS_36_wea(D2PHIDn1),
      AS_D2PHIDin_writeaddr => AS_36_writeaddr(D2PHIDn1),
      AS_D2PHIDin_din       => AS_36_din(D2PHIDn1),
      AS_D3PHIAin_wea       => AS_36_wea(D3PHIAn1),
      AS_D3PHIAin_writeaddr => AS_36_writeaddr(D3PHIAn1),
      AS_D3PHIAin_din       => AS_36_din(D3PHIAn1),
      AS_D3PHIBin_wea       => AS_36_wea(D3PHIBn1),
      AS_D3PHIBin_writeaddr => AS_36_writeaddr(D3PHIBn1),
      AS_D3PHIBin_din       => AS_36_din(D3PHIBn1),
      AS_D3PHICin_wea       => AS_36_wea(D3PHICn1),
      AS_D3PHICin_writeaddr => AS_36_writeaddr(D3PHICn1),
      AS_D3PHICin_din       => AS_36_din(D3PHICn1),
      AS_D3PHIDin_wea       => AS_36_wea(D3PHIDn1),
      AS_D3PHIDin_writeaddr => AS_36_writeaddr(D3PHIDn1),
      AS_D3PHIDin_din       => AS_36_din(D3PHIDn1),
      AS_D4PHIAin_wea       => AS_36_wea(D4PHIAn1),
      AS_D4PHIAin_writeaddr => AS_36_writeaddr(D4PHIAn1),
      AS_D4PHIAin_din       => AS_36_din(D4PHIAn1),
      AS_D4PHIBin_wea       => AS_36_wea(D4PHIBn1),
      AS_D4PHIBin_writeaddr => AS_36_writeaddr(D4PHIBn1),
      AS_D4PHIBin_din       => AS_36_din(D4PHIBn1),
      AS_D4PHICin_wea       => AS_36_wea(D4PHICn1),
      AS_D4PHICin_writeaddr => AS_36_writeaddr(D4PHICn1),
      AS_D4PHICin_din       => AS_36_din(D4PHICn1),
      AS_D4PHIDin_wea       => AS_36_wea(D4PHIDn1),
      AS_D4PHIDin_writeaddr => AS_36_writeaddr(D4PHIDn1),
      AS_D4PHIDin_din       => AS_36_din(D4PHIDn1),
      AS_D5PHIAin_wea       => AS_36_wea(D5PHIAn1),
      AS_D5PHIAin_writeaddr => AS_36_writeaddr(D5PHIAn1),
      AS_D5PHIAin_din       => AS_36_din(D5PHIAn1),
      AS_D5PHIBin_wea       => AS_36_wea(D5PHIBn1),
      AS_D5PHIBin_writeaddr => AS_36_writeaddr(D5PHIBn1),
      AS_D5PHIBin_din       => AS_36_din(D5PHIBn1),
      AS_D5PHICin_wea       => AS_36_wea(D5PHICn1),
      AS_D5PHICin_writeaddr => AS_36_writeaddr(D5PHICn1),
      AS_D5PHICin_din       => AS_36_din(D5PHICn1),
      AS_D5PHIDin_wea       => AS_36_wea(D5PHIDn1),
      AS_D5PHIDin_writeaddr => AS_36_writeaddr(D5PHIDn1),
      AS_D5PHIDin_din       => AS_36_din(D5PHIDn1),
      MPAR_L1L2ABCin_wea        => MPAR_73_wea(L1L2ABC),
      MPAR_L1L2ABCin_writeaddr  => MPAR_73_writeaddr(L1L2ABC),
      MPAR_L1L2ABCin_din        => MPAR_73_din(L1L2ABC),
      MPAR_L1L2DEin_wea         => MPAR_73_wea(L1L2DE),
      MPAR_L1L2DEin_writeaddr   => MPAR_73_writeaddr(L1L2DE),
      MPAR_L1L2DEin_din         => MPAR_73_din(L1L2DE),
      MPAR_L1L2Fin_wea          => MPAR_73_wea(L1L2F),
      MPAR_L1L2Fin_writeaddr    => MPAR_73_writeaddr(L1L2F),
      MPAR_L1L2Fin_din          => MPAR_73_din(L1L2F),
      MPAR_L1L2Gin_wea          => MPAR_73_wea(L1L2G),
      MPAR_L1L2Gin_writeaddr    => MPAR_73_writeaddr(L1L2G),
      MPAR_L1L2Gin_din          => MPAR_73_din(L1L2G),
      MPAR_L1L2HIin_wea         => MPAR_73_wea(L1L2HI),
      MPAR_L1L2HIin_writeaddr   => MPAR_73_writeaddr(L1L2HI),
      MPAR_L1L2HIin_din         => MPAR_73_din(L1L2HI),
      MPAR_L1L2JKLin_wea        => MPAR_73_wea(L1L2JKL),
      MPAR_L1L2JKLin_writeaddr  => MPAR_73_writeaddr(L1L2JKL),
      MPAR_L1L2JKLin_din        => MPAR_73_din(L1L2JKL),
      MPAR_L2L3ABCDin_wea       => MPAR_73_wea(L2L3ABCD),
      MPAR_L2L3ABCDin_writeaddr => MPAR_73_writeaddr(L2L3ABCD),
      MPAR_L2L3ABCDin_din       => MPAR_73_din(L2L3ABCD),
      MPAR_L3L4ABin_wea         => MPAR_73_wea(L3L4AB),
      MPAR_L3L4ABin_writeaddr   => MPAR_73_writeaddr(L3L4AB),
      MPAR_L3L4ABin_din         => MPAR_73_din(L3L4AB),
      MPAR_L3L4CDin_wea         => MPAR_73_wea(L3L4CD),
      MPAR_L3L4CDin_writeaddr   => MPAR_73_writeaddr(L3L4CD),
      MPAR_L3L4CDin_din         => MPAR_73_din(L3L4CD),
      MPAR_L5L6ABCDin_wea       => MPAR_73_wea(L5L6ABCD),
      MPAR_L5L6ABCDin_writeaddr => MPAR_73_writeaddr(L5L6ABCD),
      MPAR_L5L6ABCDin_din       => MPAR_73_din(L5L6ABCD),
      MPAR_D1D2ABCDin_wea       => MPAR_73_wea(D1D2ABCD),
      MPAR_D1D2ABCDin_writeaddr => MPAR_73_writeaddr(D1D2ABCD),
      MPAR_D1D2ABCDin_din       => MPAR_73_din(D1D2ABCD),
      MPAR_D3D4ABCDin_wea       => MPAR_73_wea(D3D4ABCD),
      MPAR_D3D4ABCDin_writeaddr => MPAR_73_writeaddr(D3D4ABCD),
      MPAR_D3D4ABCDin_din       => MPAR_73_din(D3D4ABCD),
      MPAR_L1D1ABCDin_wea       => MPAR_73_wea(L1D1ABCD),
      MPAR_L1D1ABCDin_writeaddr => MPAR_73_writeaddr(L1D1ABCD),
      MPAR_L1D1ABCDin_din       => MPAR_73_din(L1D1ABCD),
      MPAR_L1D1EFGHin_wea       => MPAR_73_wea(L1D1EFGH),
      MPAR_L1D1EFGHin_writeaddr => MPAR_73_writeaddr(L1D1EFGH),
      MPAR_L1D1EFGHin_din       => MPAR_73_din(L1D1EFGH),
      MPAR_L2D1ABCDin_wea       => MPAR_73_wea(L2D1ABCD),
      MPAR_L2D1ABCDin_writeaddr => MPAR_73_writeaddr(L2D1ABCD),
      MPAR_L2D1ABCDin_din       => MPAR_73_din(L2D1ABCD),
      TW_L1L2_stream_AV_din     => TW_104_stream_AV_din(L1L2),
      TW_L1L2_stream_A_full_neg => TW_104_stream_A_full_neg(L1L2),
      TW_L1L2_stream_A_write    => TW_104_stream_A_write(L1L2),
      TW_L2L3_stream_AV_din     => TW_104_stream_AV_din(L2L3),
      TW_L2L3_stream_A_full_neg => TW_104_stream_A_full_neg(L2L3),
      TW_L2L3_stream_A_write    => TW_104_stream_A_write(L2L3),
      TW_L3L4_stream_AV_din     => TW_104_stream_AV_din(L3L4),
      TW_L3L4_stream_A_full_neg => TW_104_stream_A_full_neg(L3L4),
      TW_L3L4_stream_A_write    => TW_104_stream_A_write(L3L4),
      TW_L5L6_stream_AV_din     => TW_104_stream_AV_din(L5L6),
      TW_L5L6_stream_A_full_neg => TW_104_stream_A_full_neg(L5L6),
      TW_L5L6_stream_A_write    => TW_104_stream_A_write(L5L6),
      TW_D1D2_stream_AV_din     => TW_104_stream_AV_din(D1D2),
      TW_D1D2_stream_A_full_neg => TW_104_stream_A_full_neg(D1D2),
      TW_D1D2_stream_A_write    => TW_104_stream_A_write(D1D2),
      TW_D3D4_stream_AV_din     => TW_104_stream_AV_din(D3D4),
      TW_D3D4_stream_A_full_neg => TW_104_stream_A_full_neg(D3D4),
      TW_D3D4_stream_A_write    => TW_104_stream_A_write(D3D4),
      TW_L1D1_stream_AV_din     => TW_104_stream_AV_din(L1D1),
      TW_L1D1_stream_A_full_neg => TW_104_stream_A_full_neg(L1D1),
      TW_L1D1_stream_A_write    => TW_104_stream_A_write(L1D1),
      TW_L2D1_stream_AV_din     => TW_104_stream_AV_din(L2D1),
      TW_L2D1_stream_A_full_neg => TW_104_stream_A_full_neg(L2D1),
      TW_L2D1_stream_A_write    => TW_104_stream_A_write(L2D1),
      DW_L1L2_D1_stream_AV_din     => DW_49_stream_AV_din(L1L2_D1),
      DW_L1L2_D1_stream_A_full_neg => DW_49_stream_A_full_neg(L1L2_D1),
      DW_L1L2_D1_stream_A_write    => DW_49_stream_A_write(L1L2_D1),
      DW_L1L2_D2_stream_AV_din     => DW_49_stream_AV_din(L1L2_D2),
      DW_L1L2_D2_stream_A_full_neg => DW_49_stream_A_full_neg(L1L2_D2),
      DW_L1L2_D2_stream_A_write    => DW_49_stream_A_write(L1L2_D2),
      DW_L1L2_D3_stream_AV_din     => DW_49_stream_AV_din(L1L2_D3),
      DW_L1L2_D3_stream_A_full_neg => DW_49_stream_A_full_neg(L1L2_D3),
      DW_L1L2_D3_stream_A_write    => DW_49_stream_A_write(L1L2_D3),
      DW_L1L2_D4_stream_AV_din     => DW_49_stream_AV_din(L1L2_D4),
      DW_L1L2_D4_stream_A_full_neg => DW_49_stream_A_full_neg(L1L2_D4),
      DW_L1L2_D4_stream_A_write    => DW_49_stream_A_write(L1L2_D4),
      DW_L2L3_D1_stream_AV_din     => DW_49_stream_AV_din(L2L3_D1),
      DW_L2L3_D1_stream_A_full_neg => DW_49_stream_A_full_neg(L2L3_D1),
      DW_L2L3_D1_stream_A_write    => DW_49_stream_A_write(L2L3_D1),
      DW_L2L3_D2_stream_AV_din     => DW_49_stream_AV_din(L2L3_D2),
      DW_L2L3_D2_stream_A_full_neg => DW_49_stream_A_full_neg(L2L3_D2),
      DW_L2L3_D2_stream_A_write    => DW_49_stream_A_write(L2L3_D2),
      DW_L2L3_D3_stream_AV_din     => DW_49_stream_AV_din(L2L3_D3),
      DW_L2L3_D3_stream_A_full_neg => DW_49_stream_A_full_neg(L2L3_D3),
      DW_L2L3_D3_stream_A_write    => DW_49_stream_A_write(L2L3_D3),
      DW_L2L3_D4_stream_AV_din     => DW_49_stream_AV_din(L2L3_D4),
      DW_L2L3_D4_stream_A_full_neg => DW_49_stream_A_full_neg(L2L3_D4),
      DW_L2L3_D4_stream_A_write    => DW_49_stream_A_write(L2L3_D4),
      DW_L3L4_D1_stream_AV_din     => DW_49_stream_AV_din(L3L4_D1),
      DW_L3L4_D1_stream_A_full_neg => DW_49_stream_A_full_neg(L3L4_D1),
      DW_L3L4_D1_stream_A_write    => DW_49_stream_A_write(L3L4_D1),
      DW_L3L4_D2_stream_AV_din     => DW_49_stream_AV_din(L3L4_D2),
      DW_L3L4_D2_stream_A_full_neg => DW_49_stream_A_full_neg(L3L4_D2),
      DW_L3L4_D2_stream_A_write    => DW_49_stream_A_write(L3L4_D2),
      DW_D1D2_D3_stream_AV_din     => DW_49_stream_AV_din(D1D2_D3),
      DW_D1D2_D3_stream_A_full_neg => DW_49_stream_A_full_neg(D1D2_D3),
      DW_D1D2_D3_stream_A_write    => DW_49_stream_A_write(D1D2_D3),
      DW_D1D2_D4_stream_AV_din     => DW_49_stream_AV_din(D1D2_D4),
      DW_D1D2_D4_stream_A_full_neg => DW_49_stream_A_full_neg(D1D2_D4),
      DW_D1D2_D4_stream_A_write    => DW_49_stream_A_write(D1D2_D4),
      DW_D1D2_D5_stream_AV_din     => DW_49_stream_AV_din(D1D2_D5),
      DW_D1D2_D5_stream_A_full_neg => DW_49_stream_A_full_neg(D1D2_D5),
      DW_D1D2_D5_stream_A_write    => DW_49_stream_A_write(D1D2_D5),
      DW_D3D4_D1_stream_AV_din     => DW_49_stream_AV_din(D3D4_D1),
      DW_D3D4_D1_stream_A_full_neg => DW_49_stream_A_full_neg(D3D4_D1),
      DW_D3D4_D1_stream_A_write    => DW_49_stream_A_write(D3D4_D1),
      DW_D3D4_D2_stream_AV_din     => DW_49_stream_AV_din(D3D4_D2),
      DW_D3D4_D2_stream_A_full_neg => DW_49_stream_A_full_neg(D3D4_D2),
      DW_D3D4_D2_stream_A_write    => DW_49_stream_A_write(D3D4_D2),
      DW_D3D4_D5_stream_AV_din     => DW_49_stream_AV_din(D3D4_D5),
      DW_D3D4_D5_stream_A_full_neg => DW_49_stream_A_full_neg(D3D4_D5),
      DW_D3D4_D5_stream_A_write    => DW_49_stream_A_write(D3D4_D5),
      DW_L1D1_D2_stream_AV_din     => DW_49_stream_AV_din(L1D1_D2),
      DW_L1D1_D2_stream_A_full_neg => DW_49_stream_A_full_neg(L1D1_D2),
      DW_L1D1_D2_stream_A_write    => DW_49_stream_A_write(L1D1_D2),
      DW_L1D1_D3_stream_AV_din     => DW_49_stream_AV_din(L1D1_D3),
      DW_L1D1_D3_stream_A_full_neg => DW_49_stream_A_full_neg(L1D1_D3),
      DW_L1D1_D3_stream_A_write    => DW_49_stream_A_write(L1D1_D3),
      DW_L1D1_D4_stream_AV_din     => DW_49_stream_AV_din(L1D1_D4),
      DW_L1D1_D4_stream_A_full_neg => DW_49_stream_A_full_neg(L1D1_D4),
      DW_L1D1_D4_stream_A_write    => DW_49_stream_A_write(L1D1_D4),
      DW_L1D1_D5_stream_AV_din     => DW_49_stream_AV_din(L1D1_D5),
      DW_L1D1_D5_stream_A_full_neg => DW_49_stream_A_full_neg(L1D1_D5),
      DW_L1D1_D5_stream_A_write    => DW_49_stream_A_write(L1D1_D5),
      DW_L2D1_D2_stream_AV_din     => DW_49_stream_AV_din(L2D1_D2),
      DW_L2D1_D2_stream_A_full_neg => DW_49_stream_A_full_neg(L2D1_D2),
      DW_L2D1_D2_stream_A_write    => DW_49_stream_A_write(L2D1_D2),
      DW_L2D1_D3_stream_AV_din     => DW_49_stream_AV_din(L2D1_D3),
      DW_L2D1_D3_stream_A_full_neg => DW_49_stream_A_full_neg(L2D1_D3),
      DW_L2D1_D3_stream_A_write    => DW_49_stream_A_write(L2D1_D3),
      DW_L2D1_D4_stream_AV_din     => DW_49_stream_AV_din(L2D1_D4),
      DW_L2D1_D4_stream_A_full_neg => DW_49_stream_A_full_neg(L2D1_D4),
      DW_L2D1_D4_stream_A_write    => DW_49_stream_A_write(L2D1_D4),
      BW_L1L2_L3_stream_AV_din     => BW_46_stream_AV_din(L1L2_L3),
      BW_L1L2_L3_stream_A_full_neg => BW_46_stream_A_full_neg(L1L2_L3),
      BW_L1L2_L3_stream_A_write    => BW_46_stream_A_write(L1L2_L3),
      BW_L1L2_L4_stream_AV_din     => BW_46_stream_AV_din(L1L2_L4),
      BW_L1L2_L4_stream_A_full_neg => BW_46_stream_A_full_neg(L1L2_L4),
      BW_L1L2_L4_stream_A_write    => BW_46_stream_A_write(L1L2_L4),
      BW_L1L2_L5_stream_AV_din     => BW_46_stream_AV_din(L1L2_L5),
      BW_L1L2_L5_stream_A_full_neg => BW_46_stream_A_full_neg(L1L2_L5),
      BW_L1L2_L5_stream_A_write    => BW_46_stream_A_write(L1L2_L5),
      BW_L1L2_L6_stream_AV_din     => BW_46_stream_AV_din(L1L2_L6),
      BW_L1L2_L6_stream_A_full_neg => BW_46_stream_A_full_neg(L1L2_L6),
      BW_L1L2_L6_stream_A_write    => BW_46_stream_A_write(L1L2_L6),
      BW_L2L3_L1_stream_AV_din     => BW_46_stream_AV_din(L2L3_L1),
      BW_L2L3_L1_stream_A_full_neg => BW_46_stream_A_full_neg(L2L3_L1),
      BW_L2L3_L1_stream_A_write    => BW_46_stream_A_write(L2L3_L1),
      BW_L2L3_L4_stream_AV_din     => BW_46_stream_AV_din(L2L3_L4),
      BW_L2L3_L4_stream_A_full_neg => BW_46_stream_A_full_neg(L2L3_L4),
      BW_L2L3_L4_stream_A_write    => BW_46_stream_A_write(L2L3_L4),
      BW_L2L3_L5_stream_AV_din     => BW_46_stream_AV_din(L2L3_L5),
      BW_L2L3_L5_stream_A_full_neg => BW_46_stream_A_full_neg(L2L3_L5),
      BW_L2L3_L5_stream_A_write    => BW_46_stream_A_write(L2L3_L5),
      BW_L3L4_L1_stream_AV_din     => BW_46_stream_AV_din(L3L4_L1),
      BW_L3L4_L1_stream_A_full_neg => BW_46_stream_A_full_neg(L3L4_L1),
      BW_L3L4_L1_stream_A_write    => BW_46_stream_A_write(L3L4_L1),
      BW_L3L4_L2_stream_AV_din     => BW_46_stream_AV_din(L3L4_L2),
      BW_L3L4_L2_stream_A_full_neg => BW_46_stream_A_full_neg(L3L4_L2),
      BW_L3L4_L2_stream_A_write    => BW_46_stream_A_write(L3L4_L2),
      BW_L3L4_L5_stream_AV_din     => BW_46_stream_AV_din(L3L4_L5),
      BW_L3L4_L5_stream_A_full_neg => BW_46_stream_A_full_neg(L3L4_L5),
      BW_L3L4_L5_stream_A_write    => BW_46_stream_A_write(L3L4_L5),
      BW_L3L4_L6_stream_AV_din     => BW_46_stream_AV_din(L3L4_L6),
      BW_L3L4_L6_stream_A_full_neg => BW_46_stream_A_full_neg(L3L4_L6),
      BW_L3L4_L6_stream_A_write    => BW_46_stream_A_write(L3L4_L6),
      BW_L5L6_L1_stream_AV_din     => BW_46_stream_AV_din(L5L6_L1),
      BW_L5L6_L1_stream_A_full_neg => BW_46_stream_A_full_neg(L5L6_L1),
      BW_L5L6_L1_stream_A_write    => BW_46_stream_A_write(L5L6_L1),
      BW_L5L6_L2_stream_AV_din     => BW_46_stream_AV_din(L5L6_L2),
      BW_L5L6_L2_stream_A_full_neg => BW_46_stream_A_full_neg(L5L6_L2),
      BW_L5L6_L2_stream_A_write    => BW_46_stream_A_write(L5L6_L2),
      BW_L5L6_L3_stream_AV_din     => BW_46_stream_AV_din(L5L6_L3),
      BW_L5L6_L3_stream_A_full_neg => BW_46_stream_A_full_neg(L5L6_L3),
      BW_L5L6_L3_stream_A_write    => BW_46_stream_A_write(L5L6_L3),
      BW_L5L6_L4_stream_AV_din     => BW_46_stream_AV_din(L5L6_L4),
      BW_L5L6_L4_stream_A_full_neg => BW_46_stream_A_full_neg(L5L6_L4),
      BW_L5L6_L4_stream_A_write    => BW_46_stream_A_write(L5L6_L4),
      BW_D1D2_L1_stream_AV_din     => BW_46_stream_AV_din(D1D2_L1),
      BW_D1D2_L1_stream_A_full_neg => BW_46_stream_A_full_neg(D1D2_L1),
      BW_D1D2_L1_stream_A_write    => BW_46_stream_A_write(D1D2_L1),
      BW_D1D2_L2_stream_AV_din     => BW_46_stream_AV_din(D1D2_L2),
      BW_D1D2_L2_stream_A_full_neg => BW_46_stream_A_full_neg(D1D2_L2),
      BW_D1D2_L2_stream_A_write    => BW_46_stream_A_write(D1D2_L2),
      BW_D3D4_L1_stream_AV_din     => BW_46_stream_AV_din(D3D4_L1),
      BW_D3D4_L1_stream_A_full_neg => BW_46_stream_A_full_neg(D3D4_L1),
      BW_D3D4_L1_stream_A_write    => BW_46_stream_A_write(D3D4_L1),
      BW_L2D1_L1_stream_AV_din     => BW_46_stream_AV_din(L2D1_L1),
      BW_L2D1_L1_stream_A_full_neg => BW_46_stream_A_full_neg(L2D1_L1),
      BW_L2D1_L1_stream_A_write    => BW_46_stream_A_write(L2D1_L1)
      );

end architecture rtl;
