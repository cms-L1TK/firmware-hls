--! Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--! User packages
use work.tf_pkg.all;
use work.memUtil_pkg.all;

entity SectorProcessor is
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    PC_start  : in std_logic;
    PC_bx_in : in std_logic_vector(2 downto 0);
    PC_bx_out : out std_logic_vector(2 downto 0);
    PC_bx_out_vld : out std_logic;
    PC_done : out std_logic;
    TB_bx_out : out std_logic_vector(2 downto 0);
    TB_bx_out_vld : out std_logic;
    TB_done   : out std_logic;
    TB_AAAA_last_track   : out std_logic;
    TB_AAAA_last_track_vld   : out std_logic;
    TB_BBBB_last_track   : out std_logic;
    TB_BBBB_last_track_vld   : out std_logic;
    AS_L1PHIAin_wea        : in t_AS_36_1b;
    AS_L1PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIAin_din       : in t_AS_36_DATA;
    AS_L1PHIBin_wea        : in t_AS_36_1b;
    AS_L1PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIBin_din       : in t_AS_36_DATA;
    AS_L1PHICin_wea        : in t_AS_36_1b;
    AS_L1PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHICin_din       : in t_AS_36_DATA;
    AS_L1PHIDin_wea        : in t_AS_36_1b;
    AS_L1PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIDin_din       : in t_AS_36_DATA;
    AS_L1PHIEin_wea        : in t_AS_36_1b;
    AS_L1PHIEin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIEin_din       : in t_AS_36_DATA;
    AS_L1PHIFin_wea        : in t_AS_36_1b;
    AS_L1PHIFin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIFin_din       : in t_AS_36_DATA;
    AS_L1PHIGin_wea        : in t_AS_36_1b;
    AS_L1PHIGin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIGin_din       : in t_AS_36_DATA;
    AS_L1PHIHin_wea        : in t_AS_36_1b;
    AS_L1PHIHin_writeaddr : in t_AS_36_ADDR;
    AS_L1PHIHin_din       : in t_AS_36_DATA;
    AS_L2PHIAin_wea        : in t_AS_36_1b;
    AS_L2PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L2PHIAin_din       : in t_AS_36_DATA;
    AS_L2PHIBin_wea        : in t_AS_36_1b;
    AS_L2PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L2PHIBin_din       : in t_AS_36_DATA;
    AS_L2PHICin_wea        : in t_AS_36_1b;
    AS_L2PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L2PHICin_din       : in t_AS_36_DATA;
    AS_L2PHIDin_wea        : in t_AS_36_1b;
    AS_L2PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L2PHIDin_din       : in t_AS_36_DATA;
    AS_L3PHIAin_wea        : in t_AS_36_1b;
    AS_L3PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L3PHIAin_din       : in t_AS_36_DATA;
    AS_L3PHIBin_wea        : in t_AS_36_1b;
    AS_L3PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L3PHIBin_din       : in t_AS_36_DATA;
    AS_L3PHICin_wea        : in t_AS_36_1b;
    AS_L3PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L3PHICin_din       : in t_AS_36_DATA;
    AS_L3PHIDin_wea        : in t_AS_36_1b;
    AS_L3PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L3PHIDin_din       : in t_AS_36_DATA;
    AS_L4PHIAin_wea        : in t_AS_36_1b;
    AS_L4PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L4PHIAin_din       : in t_AS_36_DATA;
    AS_L4PHIBin_wea        : in t_AS_36_1b;
    AS_L4PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L4PHIBin_din       : in t_AS_36_DATA;
    AS_L4PHICin_wea        : in t_AS_36_1b;
    AS_L4PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L4PHICin_din       : in t_AS_36_DATA;
    AS_L4PHIDin_wea        : in t_AS_36_1b;
    AS_L4PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L4PHIDin_din       : in t_AS_36_DATA;
    AS_L5PHIAin_wea        : in t_AS_36_1b;
    AS_L5PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L5PHIAin_din       : in t_AS_36_DATA;
    AS_L5PHIBin_wea        : in t_AS_36_1b;
    AS_L5PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L5PHIBin_din       : in t_AS_36_DATA;
    AS_L5PHICin_wea        : in t_AS_36_1b;
    AS_L5PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L5PHICin_din       : in t_AS_36_DATA;
    AS_L5PHIDin_wea        : in t_AS_36_1b;
    AS_L5PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L5PHIDin_din       : in t_AS_36_DATA;
    AS_L6PHIAin_wea        : in t_AS_36_1b;
    AS_L6PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_L6PHIAin_din       : in t_AS_36_DATA;
    AS_L6PHIBin_wea        : in t_AS_36_1b;
    AS_L6PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_L6PHIBin_din       : in t_AS_36_DATA;
    AS_L6PHICin_wea        : in t_AS_36_1b;
    AS_L6PHICin_writeaddr : in t_AS_36_ADDR;
    AS_L6PHICin_din       : in t_AS_36_DATA;
    AS_L6PHIDin_wea        : in t_AS_36_1b;
    AS_L6PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_L6PHIDin_din       : in t_AS_36_DATA;
    AS_D1PHIAin_wea        : in t_AS_36_1b;
    AS_D1PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_D1PHIAin_din       : in t_AS_36_DATA;
    AS_D1PHIBin_wea        : in t_AS_36_1b;
    AS_D1PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_D1PHIBin_din       : in t_AS_36_DATA;
    AS_D1PHICin_wea        : in t_AS_36_1b;
    AS_D1PHICin_writeaddr : in t_AS_36_ADDR;
    AS_D1PHICin_din       : in t_AS_36_DATA;
    AS_D1PHIDin_wea        : in t_AS_36_1b;
    AS_D1PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_D1PHIDin_din       : in t_AS_36_DATA;
    AS_D2PHIAin_wea        : in t_AS_36_1b;
    AS_D2PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_D2PHIAin_din       : in t_AS_36_DATA;
    AS_D2PHIBin_wea        : in t_AS_36_1b;
    AS_D2PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_D2PHIBin_din       : in t_AS_36_DATA;
    AS_D2PHICin_wea        : in t_AS_36_1b;
    AS_D2PHICin_writeaddr : in t_AS_36_ADDR;
    AS_D2PHICin_din       : in t_AS_36_DATA;
    AS_D2PHIDin_wea        : in t_AS_36_1b;
    AS_D2PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_D2PHIDin_din       : in t_AS_36_DATA;
    AS_D3PHIAin_wea        : in t_AS_36_1b;
    AS_D3PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_D3PHIAin_din       : in t_AS_36_DATA;
    AS_D3PHIBin_wea        : in t_AS_36_1b;
    AS_D3PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_D3PHIBin_din       : in t_AS_36_DATA;
    AS_D3PHICin_wea        : in t_AS_36_1b;
    AS_D3PHICin_writeaddr : in t_AS_36_ADDR;
    AS_D3PHICin_din       : in t_AS_36_DATA;
    AS_D3PHIDin_wea        : in t_AS_36_1b;
    AS_D3PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_D3PHIDin_din       : in t_AS_36_DATA;
    AS_D4PHIAin_wea        : in t_AS_36_1b;
    AS_D4PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_D4PHIAin_din       : in t_AS_36_DATA;
    AS_D4PHIBin_wea        : in t_AS_36_1b;
    AS_D4PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_D4PHIBin_din       : in t_AS_36_DATA;
    AS_D4PHICin_wea        : in t_AS_36_1b;
    AS_D4PHICin_writeaddr : in t_AS_36_ADDR;
    AS_D4PHICin_din       : in t_AS_36_DATA;
    AS_D4PHIDin_wea        : in t_AS_36_1b;
    AS_D4PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_D4PHIDin_din       : in t_AS_36_DATA;
    AS_D5PHIAin_wea        : in t_AS_36_1b;
    AS_D5PHIAin_writeaddr : in t_AS_36_ADDR;
    AS_D5PHIAin_din       : in t_AS_36_DATA;
    AS_D5PHIBin_wea        : in t_AS_36_1b;
    AS_D5PHIBin_writeaddr : in t_AS_36_ADDR;
    AS_D5PHIBin_din       : in t_AS_36_DATA;
    AS_D5PHICin_wea        : in t_AS_36_1b;
    AS_D5PHICin_writeaddr : in t_AS_36_ADDR;
    AS_D5PHICin_din       : in t_AS_36_DATA;
    AS_D5PHIDin_wea        : in t_AS_36_1b;
    AS_D5PHIDin_writeaddr : in t_AS_36_ADDR;
    AS_D5PHIDin_din       : in t_AS_36_DATA;
    MPAR_L1L2ABCin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2ABCin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2ABCin_din       : in t_MPAR_73_DATA;
    MPAR_L1L2DEin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2DEin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2DEin_din       : in t_MPAR_73_DATA;
    MPAR_L1L2Fin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2Fin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2Fin_din       : in t_MPAR_73_DATA;
    MPAR_L1L2Gin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2Gin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2Gin_din       : in t_MPAR_73_DATA;
    MPAR_L1L2HIin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2HIin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2HIin_din       : in t_MPAR_73_DATA;
    MPAR_L1L2JKLin_wea        : in t_MPAR_73_1b;
    MPAR_L1L2JKLin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1L2JKLin_din       : in t_MPAR_73_DATA;
    MPAR_L2L3ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_L2L3ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L2L3ABCDin_din       : in t_MPAR_73_DATA;
    MPAR_L3L4ABin_wea        : in t_MPAR_73_1b;
    MPAR_L3L4ABin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L3L4ABin_din       : in t_MPAR_73_DATA;
    MPAR_L3L4CDin_wea        : in t_MPAR_73_1b;
    MPAR_L3L4CDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L3L4CDin_din       : in t_MPAR_73_DATA;
    MPAR_L5L6ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_L5L6ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L5L6ABCDin_din       : in t_MPAR_73_DATA;
    MPAR_D1D2ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_D1D2ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_D1D2ABCDin_din       : in t_MPAR_73_DATA;
    MPAR_D3D4ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_D3D4ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_D3D4ABCDin_din       : in t_MPAR_73_DATA;
    MPAR_L1D1ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_L1D1ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1D1ABCDin_din       : in t_MPAR_73_DATA;
    MPAR_L1D1EFGHin_wea        : in t_MPAR_73_1b;
    MPAR_L1D1EFGHin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L1D1EFGHin_din       : in t_MPAR_73_DATA;
    MPAR_L2D1ABCDin_wea        : in t_MPAR_73_1b;
    MPAR_L2D1ABCDin_writeaddr : in t_MPAR_73_ADDR;
    MPAR_L2D1ABCDin_din       : in t_MPAR_73_DATA;
    TW_AAAA_stream_AV_din       : out t_TW_113_DATA;
    TW_AAAA_stream_A_full_neg   : in t_TW_113_1b;
    TW_AAAA_stream_A_write      : out t_TW_113_1b;
    TW_BBBB_stream_AV_din       : out t_TW_113_DATA;
    TW_BBBB_stream_A_full_neg   : in t_TW_113_1b;
    TW_BBBB_stream_A_write      : out t_TW_113_1b;
    DW_AAAA_D1_stream_AV_din       : out t_DW_49_DATA;
    DW_AAAA_D1_stream_A_full_neg   : in t_DW_49_1b;
    DW_AAAA_D1_stream_A_write      : out t_DW_49_1b;
    DW_AAAA_D2_stream_AV_din       : out t_DW_49_DATA;
    DW_AAAA_D2_stream_A_full_neg   : in t_DW_49_1b;
    DW_AAAA_D2_stream_A_write      : out t_DW_49_1b;
    DW_AAAA_D3_stream_AV_din       : out t_DW_49_DATA;
    DW_AAAA_D3_stream_A_full_neg   : in t_DW_49_1b;
    DW_AAAA_D3_stream_A_write      : out t_DW_49_1b;
    DW_AAAA_D4_stream_AV_din       : out t_DW_49_DATA;
    DW_AAAA_D4_stream_A_full_neg   : in t_DW_49_1b;
    DW_AAAA_D4_stream_A_write      : out t_DW_49_1b;
    DW_AAAA_D5_stream_AV_din       : out t_DW_49_DATA;
    DW_AAAA_D5_stream_A_full_neg   : in t_DW_49_1b;
    DW_AAAA_D5_stream_A_write      : out t_DW_49_1b;
    DW_BBBB_D1_stream_AV_din       : out t_DW_49_DATA;
    DW_BBBB_D1_stream_A_full_neg   : in t_DW_49_1b;
    DW_BBBB_D1_stream_A_write      : out t_DW_49_1b;
    DW_BBBB_D2_stream_AV_din       : out t_DW_49_DATA;
    DW_BBBB_D2_stream_A_full_neg   : in t_DW_49_1b;
    DW_BBBB_D2_stream_A_write      : out t_DW_49_1b;
    DW_BBBB_D3_stream_AV_din       : out t_DW_49_DATA;
    DW_BBBB_D3_stream_A_full_neg   : in t_DW_49_1b;
    DW_BBBB_D3_stream_A_write      : out t_DW_49_1b;
    DW_BBBB_D4_stream_AV_din       : out t_DW_49_DATA;
    DW_BBBB_D4_stream_A_full_neg   : in t_DW_49_1b;
    DW_BBBB_D4_stream_A_write      : out t_DW_49_1b;
    DW_BBBB_D5_stream_AV_din       : out t_DW_49_DATA;
    DW_BBBB_D5_stream_A_full_neg   : in t_DW_49_1b;
    DW_BBBB_D5_stream_A_write      : out t_DW_49_1b;
    BW_AAAA_L1_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L1_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L1_stream_A_write      : out t_BW_46_1b;
    BW_AAAA_L2_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L2_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L2_stream_A_write      : out t_BW_46_1b;
    BW_AAAA_L3_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L3_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L3_stream_A_write      : out t_BW_46_1b;
    BW_AAAA_L4_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L4_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L4_stream_A_write      : out t_BW_46_1b;
    BW_AAAA_L5_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L5_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L5_stream_A_write      : out t_BW_46_1b;
    BW_AAAA_L6_stream_AV_din       : out t_BW_46_DATA;
    BW_AAAA_L6_stream_A_full_neg   : in t_BW_46_1b;
    BW_AAAA_L6_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L1_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L1_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L1_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L2_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L2_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L2_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L3_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L3_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L3_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L4_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L4_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L4_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L5_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L5_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L5_stream_A_write      : out t_BW_46_1b;
    BW_BBBB_L6_stream_AV_din       : out t_BW_46_DATA;
    BW_BBBB_L6_stream_A_full_neg   : in t_BW_46_1b;
    BW_BBBB_L6_stream_A_write      : out t_BW_46_1b
  );
end SectorProcessor;

architecture rtl of SectorProcessor is

  signal AS_L1PHIAin_start                   : std_logic;
  signal AS_L1PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIAin_valid        : STD_LOGIC;
  signal AS_L1PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIBin_start                   : std_logic;
  signal AS_L1PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIBin_valid        : STD_LOGIC;
  signal AS_L1PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHICin_start                   : std_logic;
  signal AS_L1PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHICin_V_as        : t_AS_36_DATA;
  signal AS_L1PHICin_valid        : STD_LOGIC;
  signal AS_L1PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIDin_start                   : std_logic;
  signal AS_L1PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIDin_valid        : STD_LOGIC;
  signal AS_L1PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIEin_start                   : std_logic;
  signal AS_L1PHIEin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIEin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIEin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIEin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIEin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIEin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIEin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIEin_valid        : STD_LOGIC;
  signal AS_L1PHIEin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIEin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIFin_start                   : std_logic;
  signal AS_L1PHIFin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIFin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIFin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIFin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIFin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIFin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIFin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIFin_valid        : STD_LOGIC;
  signal AS_L1PHIFin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIFin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIGin_start                   : std_logic;
  signal AS_L1PHIGin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIGin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIGin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIGin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIGin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIGin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIGin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIGin_valid        : STD_LOGIC;
  signal AS_L1PHIGin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIGin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIHin_start                   : std_logic;
  signal AS_L1PHIHin_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIHin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIHin_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIHin_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIHin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIHin_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIHin_V_as        : t_AS_36_DATA;
  signal AS_L1PHIHin_valid        : STD_LOGIC;
  signal AS_L1PHIHin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L1PHIHin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIAin_start                   : std_logic;
  signal AS_L2PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L2PHIAin_valid        : STD_LOGIC;
  signal AS_L2PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L2PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIBin_start                   : std_logic;
  signal AS_L2PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L2PHIBin_valid        : STD_LOGIC;
  signal AS_L2PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L2PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHICin_start                   : std_logic;
  signal AS_L2PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L2PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L2PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L2PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L2PHICin_V_as        : t_AS_36_DATA;
  signal AS_L2PHICin_valid        : STD_LOGIC;
  signal AS_L2PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L2PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIDin_start                   : std_logic;
  signal AS_L2PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L2PHIDin_valid        : STD_LOGIC;
  signal AS_L2PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L2PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIAin_start                   : std_logic;
  signal AS_L3PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L3PHIAin_valid        : STD_LOGIC;
  signal AS_L3PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L3PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIBin_start                   : std_logic;
  signal AS_L3PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L3PHIBin_valid        : STD_LOGIC;
  signal AS_L3PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L3PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHICin_start                   : std_logic;
  signal AS_L3PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L3PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L3PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L3PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L3PHICin_V_as        : t_AS_36_DATA;
  signal AS_L3PHICin_valid        : STD_LOGIC;
  signal AS_L3PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L3PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIDin_start                   : std_logic;
  signal AS_L3PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L3PHIDin_valid        : STD_LOGIC;
  signal AS_L3PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L3PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIAin_start                   : std_logic;
  signal AS_L4PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L4PHIAin_valid        : STD_LOGIC;
  signal AS_L4PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L4PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIBin_start                   : std_logic;
  signal AS_L4PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L4PHIBin_valid        : STD_LOGIC;
  signal AS_L4PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L4PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHICin_start                   : std_logic;
  signal AS_L4PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L4PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L4PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L4PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L4PHICin_V_as        : t_AS_36_DATA;
  signal AS_L4PHICin_valid        : STD_LOGIC;
  signal AS_L4PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L4PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIDin_start                   : std_logic;
  signal AS_L4PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L4PHIDin_valid        : STD_LOGIC;
  signal AS_L4PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L4PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIAin_start                   : std_logic;
  signal AS_L5PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L5PHIAin_valid        : STD_LOGIC;
  signal AS_L5PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L5PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIBin_start                   : std_logic;
  signal AS_L5PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L5PHIBin_valid        : STD_LOGIC;
  signal AS_L5PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L5PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHICin_start                   : std_logic;
  signal AS_L5PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L5PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L5PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L5PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L5PHICin_V_as        : t_AS_36_DATA;
  signal AS_L5PHICin_valid        : STD_LOGIC;
  signal AS_L5PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L5PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIDin_start                   : std_logic;
  signal AS_L5PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L5PHIDin_valid        : STD_LOGIC;
  signal AS_L5PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L5PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIAin_start                   : std_logic;
  signal AS_L6PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIAin_V_as        : t_AS_36_DATA;
  signal AS_L6PHIAin_valid        : STD_LOGIC;
  signal AS_L6PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L6PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIBin_start                   : std_logic;
  signal AS_L6PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIBin_V_as        : t_AS_36_DATA;
  signal AS_L6PHIBin_valid        : STD_LOGIC;
  signal AS_L6PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L6PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHICin_start                   : std_logic;
  signal AS_L6PHICin_wea_delay          : t_AS_36_1b;
  signal AS_L6PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHICin_din_delay         : t_AS_36_DATA;
  signal AS_L6PHICin_enb          : t_AS_36_1b := '1';
  signal AS_L6PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHICin_V_dout        : t_AS_36_DATA;
  signal AS_L6PHICin_V_as        : t_AS_36_DATA;
  signal AS_L6PHICin_valid        : STD_LOGIC;
  signal AS_L6PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L6PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIDin_start                   : std_logic;
  signal AS_L6PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIDin_V_as        : t_AS_36_DATA;
  signal AS_L6PHIDin_valid        : STD_LOGIC;
  signal AS_L6PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_L6PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIAin_start                   : std_logic;
  signal AS_D1PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIAin_V_as        : t_AS_36_DATA;
  signal AS_D1PHIAin_valid        : STD_LOGIC;
  signal AS_D1PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D1PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIBin_start                   : std_logic;
  signal AS_D1PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIBin_V_as        : t_AS_36_DATA;
  signal AS_D1PHIBin_valid        : STD_LOGIC;
  signal AS_D1PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D1PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHICin_start                   : std_logic;
  signal AS_D1PHICin_wea_delay          : t_AS_36_1b;
  signal AS_D1PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHICin_din_delay         : t_AS_36_DATA;
  signal AS_D1PHICin_enb          : t_AS_36_1b := '1';
  signal AS_D1PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHICin_V_dout        : t_AS_36_DATA;
  signal AS_D1PHICin_V_as        : t_AS_36_DATA;
  signal AS_D1PHICin_valid        : STD_LOGIC;
  signal AS_D1PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D1PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIDin_start                   : std_logic;
  signal AS_D1PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIDin_V_as        : t_AS_36_DATA;
  signal AS_D1PHIDin_valid        : STD_LOGIC;
  signal AS_D1PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D1PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIAin_start                   : std_logic;
  signal AS_D2PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIAin_V_as        : t_AS_36_DATA;
  signal AS_D2PHIAin_valid        : STD_LOGIC;
  signal AS_D2PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D2PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIBin_start                   : std_logic;
  signal AS_D2PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIBin_V_as        : t_AS_36_DATA;
  signal AS_D2PHIBin_valid        : STD_LOGIC;
  signal AS_D2PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D2PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHICin_start                   : std_logic;
  signal AS_D2PHICin_wea_delay          : t_AS_36_1b;
  signal AS_D2PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHICin_din_delay         : t_AS_36_DATA;
  signal AS_D2PHICin_enb          : t_AS_36_1b := '1';
  signal AS_D2PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHICin_V_dout        : t_AS_36_DATA;
  signal AS_D2PHICin_V_as        : t_AS_36_DATA;
  signal AS_D2PHICin_valid        : STD_LOGIC;
  signal AS_D2PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D2PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIDin_start                   : std_logic;
  signal AS_D2PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIDin_V_as        : t_AS_36_DATA;
  signal AS_D2PHIDin_valid        : STD_LOGIC;
  signal AS_D2PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D2PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIAin_start                   : std_logic;
  signal AS_D3PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIAin_V_as        : t_AS_36_DATA;
  signal AS_D3PHIAin_valid        : STD_LOGIC;
  signal AS_D3PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D3PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIBin_start                   : std_logic;
  signal AS_D3PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIBin_V_as        : t_AS_36_DATA;
  signal AS_D3PHIBin_valid        : STD_LOGIC;
  signal AS_D3PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D3PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHICin_start                   : std_logic;
  signal AS_D3PHICin_wea_delay          : t_AS_36_1b;
  signal AS_D3PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHICin_din_delay         : t_AS_36_DATA;
  signal AS_D3PHICin_enb          : t_AS_36_1b := '1';
  signal AS_D3PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHICin_V_dout        : t_AS_36_DATA;
  signal AS_D3PHICin_V_as        : t_AS_36_DATA;
  signal AS_D3PHICin_valid        : STD_LOGIC;
  signal AS_D3PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D3PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIDin_start                   : std_logic;
  signal AS_D3PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIDin_V_as        : t_AS_36_DATA;
  signal AS_D3PHIDin_valid        : STD_LOGIC;
  signal AS_D3PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D3PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIAin_start                   : std_logic;
  signal AS_D4PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIAin_V_as        : t_AS_36_DATA;
  signal AS_D4PHIAin_valid        : STD_LOGIC;
  signal AS_D4PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D4PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIBin_start                   : std_logic;
  signal AS_D4PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIBin_V_as        : t_AS_36_DATA;
  signal AS_D4PHIBin_valid        : STD_LOGIC;
  signal AS_D4PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D4PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHICin_start                   : std_logic;
  signal AS_D4PHICin_wea_delay          : t_AS_36_1b;
  signal AS_D4PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHICin_din_delay         : t_AS_36_DATA;
  signal AS_D4PHICin_enb          : t_AS_36_1b := '1';
  signal AS_D4PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHICin_V_dout        : t_AS_36_DATA;
  signal AS_D4PHICin_V_as        : t_AS_36_DATA;
  signal AS_D4PHICin_valid        : STD_LOGIC;
  signal AS_D4PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D4PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIDin_start                   : std_logic;
  signal AS_D4PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIDin_V_as        : t_AS_36_DATA;
  signal AS_D4PHIDin_valid        : STD_LOGIC;
  signal AS_D4PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D4PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIAin_start                   : std_logic;
  signal AS_D5PHIAin_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIAin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIAin_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIAin_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIAin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIAin_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIAin_V_as        : t_AS_36_DATA;
  signal AS_D5PHIAin_valid        : STD_LOGIC;
  signal AS_D5PHIAin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D5PHIAin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIBin_start                   : std_logic;
  signal AS_D5PHIBin_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIBin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIBin_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIBin_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIBin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIBin_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIBin_V_as        : t_AS_36_DATA;
  signal AS_D5PHIBin_valid        : STD_LOGIC;
  signal AS_D5PHIBin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D5PHIBin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHICin_start                   : std_logic;
  signal AS_D5PHICin_wea_delay          : t_AS_36_1b;
  signal AS_D5PHICin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHICin_din_delay         : t_AS_36_DATA;
  signal AS_D5PHICin_enb          : t_AS_36_1b := '1';
  signal AS_D5PHICin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHICin_V_dout        : t_AS_36_DATA;
  signal AS_D5PHICin_V_as        : t_AS_36_DATA;
  signal AS_D5PHICin_valid        : STD_LOGIC;
  signal AS_D5PHICin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D5PHICin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIDin_start                   : std_logic;
  signal AS_D5PHIDin_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIDin_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIDin_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIDin_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIDin_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIDin_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIDin_V_as        : t_AS_36_DATA;
  signal AS_D5PHIDin_valid        : STD_LOGIC;
  signal AS_D5PHIDin_index        : STD_LOGIC_VECTOR(31 downto 0);
  signal AS_D5PHIDin_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIAn2_start                   : std_logic;
  signal AS_L1PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIAn2_wea          : t_AS_36_1b;
  signal AS_L1PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIAn2_din         : t_AS_36_DATA;
  signal AS_L1PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIBn2_start                   : std_logic;
  signal AS_L1PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIBn2_wea          : t_AS_36_1b;
  signal AS_L1PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIBn2_din         : t_AS_36_DATA;
  signal AS_L1PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHICn2_start                   : std_logic;
  signal AS_L1PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHICn2_wea          : t_AS_36_1b;
  signal AS_L1PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHICn2_din         : t_AS_36_DATA;
  signal AS_L1PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIDn2_start                   : std_logic;
  signal AS_L1PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIDn2_wea          : t_AS_36_1b;
  signal AS_L1PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIDn2_din         : t_AS_36_DATA;
  signal AS_L1PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIEn2_start                   : std_logic;
  signal AS_L1PHIEn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIEn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIEn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIEn2_wea          : t_AS_36_1b;
  signal AS_L1PHIEn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIEn2_din         : t_AS_36_DATA;
  signal AS_L1PHIEn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIEn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIEn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIEn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIFn2_start                   : std_logic;
  signal AS_L1PHIFn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIFn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIFn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIFn2_wea          : t_AS_36_1b;
  signal AS_L1PHIFn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIFn2_din         : t_AS_36_DATA;
  signal AS_L1PHIFn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIFn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIFn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIFn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIGn2_start                   : std_logic;
  signal AS_L1PHIGn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIGn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIGn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIGn2_wea          : t_AS_36_1b;
  signal AS_L1PHIGn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIGn2_din         : t_AS_36_DATA;
  signal AS_L1PHIGn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIGn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIGn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIGn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIHn2_start                   : std_logic;
  signal AS_L1PHIHn2_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIHn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIHn2_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIHn2_wea          : t_AS_36_1b;
  signal AS_L1PHIHn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIHn2_din         : t_AS_36_DATA;
  signal AS_L1PHIHn2_enb          : t_AS_36_1b := '1';
  signal AS_L1PHIHn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L1PHIHn2_V_dout        : t_AS_36_DATA;
  signal AS_L1PHIHn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIAn2_start                   : std_logic;
  signal AS_L2PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIAn2_wea          : t_AS_36_1b;
  signal AS_L2PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIAn2_din         : t_AS_36_DATA;
  signal AS_L2PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIBn2_start                   : std_logic;
  signal AS_L2PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIBn2_wea          : t_AS_36_1b;
  signal AS_L2PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIBn2_din         : t_AS_36_DATA;
  signal AS_L2PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHICn2_start                   : std_logic;
  signal AS_L2PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L2PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L2PHICn2_wea          : t_AS_36_1b;
  signal AS_L2PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHICn2_din         : t_AS_36_DATA;
  signal AS_L2PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L2PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L2PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIDn2_start                   : std_logic;
  signal AS_L2PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIDn2_wea          : t_AS_36_1b;
  signal AS_L2PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIDn2_din         : t_AS_36_DATA;
  signal AS_L2PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIAn2_start                   : std_logic;
  signal AS_L3PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIAn2_wea          : t_AS_36_1b;
  signal AS_L3PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIAn2_din         : t_AS_36_DATA;
  signal AS_L3PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIBn2_start                   : std_logic;
  signal AS_L3PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIBn2_wea          : t_AS_36_1b;
  signal AS_L3PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIBn2_din         : t_AS_36_DATA;
  signal AS_L3PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHICn2_start                   : std_logic;
  signal AS_L3PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L3PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L3PHICn2_wea          : t_AS_36_1b;
  signal AS_L3PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHICn2_din         : t_AS_36_DATA;
  signal AS_L3PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L3PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L3PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIDn2_start                   : std_logic;
  signal AS_L3PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIDn2_wea          : t_AS_36_1b;
  signal AS_L3PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIDn2_din         : t_AS_36_DATA;
  signal AS_L3PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIAn2_start                   : std_logic;
  signal AS_L4PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIAn2_wea          : t_AS_36_1b;
  signal AS_L4PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIAn2_din         : t_AS_36_DATA;
  signal AS_L4PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIBn2_start                   : std_logic;
  signal AS_L4PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIBn2_wea          : t_AS_36_1b;
  signal AS_L4PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIBn2_din         : t_AS_36_DATA;
  signal AS_L4PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHICn2_start                   : std_logic;
  signal AS_L4PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L4PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L4PHICn2_wea          : t_AS_36_1b;
  signal AS_L4PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHICn2_din         : t_AS_36_DATA;
  signal AS_L4PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L4PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L4PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIDn2_start                   : std_logic;
  signal AS_L4PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIDn2_wea          : t_AS_36_1b;
  signal AS_L4PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIDn2_din         : t_AS_36_DATA;
  signal AS_L4PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIAn2_start                   : std_logic;
  signal AS_L5PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIAn2_wea          : t_AS_36_1b;
  signal AS_L5PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIAn2_din         : t_AS_36_DATA;
  signal AS_L5PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIBn2_start                   : std_logic;
  signal AS_L5PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIBn2_wea          : t_AS_36_1b;
  signal AS_L5PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIBn2_din         : t_AS_36_DATA;
  signal AS_L5PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHICn2_start                   : std_logic;
  signal AS_L5PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L5PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L5PHICn2_wea          : t_AS_36_1b;
  signal AS_L5PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHICn2_din         : t_AS_36_DATA;
  signal AS_L5PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L5PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L5PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIDn2_start                   : std_logic;
  signal AS_L5PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIDn2_wea          : t_AS_36_1b;
  signal AS_L5PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIDn2_din         : t_AS_36_DATA;
  signal AS_L5PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L5PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L5PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L5PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIAn2_start                   : std_logic;
  signal AS_L6PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIAn2_wea          : t_AS_36_1b;
  signal AS_L6PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIAn2_din         : t_AS_36_DATA;
  signal AS_L6PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIBn2_start                   : std_logic;
  signal AS_L6PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIBn2_wea          : t_AS_36_1b;
  signal AS_L6PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIBn2_din         : t_AS_36_DATA;
  signal AS_L6PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHICn2_start                   : std_logic;
  signal AS_L6PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_L6PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_L6PHICn2_wea          : t_AS_36_1b;
  signal AS_L6PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHICn2_din         : t_AS_36_DATA;
  signal AS_L6PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_L6PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_L6PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIDn2_start                   : std_logic;
  signal AS_L6PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIDn2_wea          : t_AS_36_1b;
  signal AS_L6PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIDn2_din         : t_AS_36_DATA;
  signal AS_L6PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIAn2_start                   : std_logic;
  signal AS_D1PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIAn2_wea          : t_AS_36_1b;
  signal AS_D1PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIAn2_din         : t_AS_36_DATA;
  signal AS_D1PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIBn2_start                   : std_logic;
  signal AS_D1PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIBn2_wea          : t_AS_36_1b;
  signal AS_D1PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIBn2_din         : t_AS_36_DATA;
  signal AS_D1PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHICn2_start                   : std_logic;
  signal AS_D1PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_D1PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_D1PHICn2_wea          : t_AS_36_1b;
  signal AS_D1PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHICn2_din         : t_AS_36_DATA;
  signal AS_D1PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_D1PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_D1PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIDn2_start                   : std_logic;
  signal AS_D1PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIDn2_wea          : t_AS_36_1b;
  signal AS_D1PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIDn2_din         : t_AS_36_DATA;
  signal AS_D1PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIAn2_start                   : std_logic;
  signal AS_D2PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIAn2_wea          : t_AS_36_1b;
  signal AS_D2PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIAn2_din         : t_AS_36_DATA;
  signal AS_D2PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIBn2_start                   : std_logic;
  signal AS_D2PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIBn2_wea          : t_AS_36_1b;
  signal AS_D2PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIBn2_din         : t_AS_36_DATA;
  signal AS_D2PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHICn2_start                   : std_logic;
  signal AS_D2PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_D2PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_D2PHICn2_wea          : t_AS_36_1b;
  signal AS_D2PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHICn2_din         : t_AS_36_DATA;
  signal AS_D2PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_D2PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_D2PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIDn2_start                   : std_logic;
  signal AS_D2PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIDn2_wea          : t_AS_36_1b;
  signal AS_D2PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIDn2_din         : t_AS_36_DATA;
  signal AS_D2PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIAn2_start                   : std_logic;
  signal AS_D3PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIAn2_wea          : t_AS_36_1b;
  signal AS_D3PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIAn2_din         : t_AS_36_DATA;
  signal AS_D3PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIBn2_start                   : std_logic;
  signal AS_D3PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIBn2_wea          : t_AS_36_1b;
  signal AS_D3PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIBn2_din         : t_AS_36_DATA;
  signal AS_D3PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHICn2_start                   : std_logic;
  signal AS_D3PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_D3PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_D3PHICn2_wea          : t_AS_36_1b;
  signal AS_D3PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHICn2_din         : t_AS_36_DATA;
  signal AS_D3PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_D3PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_D3PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIDn2_start                   : std_logic;
  signal AS_D3PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIDn2_wea          : t_AS_36_1b;
  signal AS_D3PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIDn2_din         : t_AS_36_DATA;
  signal AS_D3PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_D3PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D3PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_D3PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIAn2_start                   : std_logic;
  signal AS_D4PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIAn2_wea          : t_AS_36_1b;
  signal AS_D4PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIAn2_din         : t_AS_36_DATA;
  signal AS_D4PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIBn2_start                   : std_logic;
  signal AS_D4PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIBn2_wea          : t_AS_36_1b;
  signal AS_D4PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIBn2_din         : t_AS_36_DATA;
  signal AS_D4PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHICn2_start                   : std_logic;
  signal AS_D4PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_D4PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_D4PHICn2_wea          : t_AS_36_1b;
  signal AS_D4PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHICn2_din         : t_AS_36_DATA;
  signal AS_D4PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_D4PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_D4PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIDn2_start                   : std_logic;
  signal AS_D4PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIDn2_wea          : t_AS_36_1b;
  signal AS_D4PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIDn2_din         : t_AS_36_DATA;
  signal AS_D4PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIAn2_start                   : std_logic;
  signal AS_D5PHIAn2_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIAn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIAn2_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIAn2_wea          : t_AS_36_1b;
  signal AS_D5PHIAn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIAn2_din         : t_AS_36_DATA;
  signal AS_D5PHIAn2_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIAn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIAn2_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIAn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIBn2_start                   : std_logic;
  signal AS_D5PHIBn2_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIBn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIBn2_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIBn2_wea          : t_AS_36_1b;
  signal AS_D5PHIBn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIBn2_din         : t_AS_36_DATA;
  signal AS_D5PHIBn2_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIBn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIBn2_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIBn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHICn2_start                   : std_logic;
  signal AS_D5PHICn2_wea_delay          : t_AS_36_1b;
  signal AS_D5PHICn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHICn2_din_delay         : t_AS_36_DATA;
  signal AS_D5PHICn2_wea          : t_AS_36_1b;
  signal AS_D5PHICn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHICn2_din         : t_AS_36_DATA;
  signal AS_D5PHICn2_enb          : t_AS_36_1b := '1';
  signal AS_D5PHICn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHICn2_V_dout        : t_AS_36_DATA;
  signal AS_D5PHICn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIDn2_start                   : std_logic;
  signal AS_D5PHIDn2_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIDn2_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIDn2_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIDn2_wea          : t_AS_36_1b;
  signal AS_D5PHIDn2_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIDn2_din         : t_AS_36_DATA;
  signal AS_D5PHIDn2_enb          : t_AS_36_1b := '1';
  signal AS_D5PHIDn2_V_readaddr    : t_AS_36_ADDR;
  signal AS_D5PHIDn2_V_dout        : t_AS_36_DATA;
  signal AS_D5PHIDn2_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal VMSME_L1PHIAn2_start                   : std_logic;
  signal VMSME_L1PHIAn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIAn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIAn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIAn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIAn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIAn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIAn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIAn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIAn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIAn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIAn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIAn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIAn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIAn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIAn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIAn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIAn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIAn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIAn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIAn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIAn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIBn2_start                   : std_logic;
  signal VMSME_L1PHIBn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIBn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIBn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIBn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIBn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIBn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIBn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIBn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIBn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIBn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIBn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIBn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIBn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIBn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIBn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIBn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIBn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIBn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIBn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIBn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIBn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHICn2_start                   : std_logic;
  signal VMSME_L1PHICn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHICn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHICn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHICn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHICn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHICn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHICn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHICn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHICn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHICn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHICn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHICn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHICn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHICn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHICn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHICn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHICn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHICn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHICn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHICn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHICn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIDn2_start                   : std_logic;
  signal VMSME_L1PHIDn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIDn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIDn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIDn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIDn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIDn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIDn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIDn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIDn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIDn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIDn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIDn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIDn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIDn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIDn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIDn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIDn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIDn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIDn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIDn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIDn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIEn2_start                   : std_logic;
  signal VMSME_L1PHIEn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIEn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIEn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIEn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIEn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIEn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIEn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIEn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIEn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIEn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIEn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIEn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIEn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIEn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIEn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIEn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIEn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIEn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIEn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIEn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIEn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIFn2_start                   : std_logic;
  signal VMSME_L1PHIFn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIFn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIFn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIFn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIFn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIFn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIFn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIFn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIFn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIFn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIFn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIFn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIFn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIFn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIFn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIFn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIFn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIFn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIFn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIFn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIFn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIGn2_start                   : std_logic;
  signal VMSME_L1PHIGn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIGn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIGn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIGn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIGn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIGn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIGn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIGn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIGn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIGn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIGn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIGn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIGn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIGn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIGn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIGn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIGn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIGn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIGn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIGn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIGn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L1PHIHn2_start                   : std_logic;
  signal VMSME_L1PHIHn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L1PHIHn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIHn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L1PHIHn2_wea          : t_VMSME_16_1b;
  signal VMSME_L1PHIHn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L1PHIHn2_din         : t_VMSME_16_DATA;
  signal VMSME_L1PHIHn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L1PHIHn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L1PHIHn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L1PHIHn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L1PHIHn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L1PHIHn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L1PHIHn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L1PHIHn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L1PHIHn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L1PHIHn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIHn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIHn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L1PHIHn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L1PHIHn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L1PHIHn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L2PHIAn2_start                   : std_logic;
  signal VMSME_L2PHIAn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L2PHIAn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIAn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L2PHIAn2_wea          : t_VMSME_16_1b;
  signal VMSME_L2PHIAn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIAn2_din         : t_VMSME_16_DATA;
  signal VMSME_L2PHIAn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L2PHIAn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L2PHIAn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L2PHIAn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L2PHIAn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L2PHIAn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L2PHIAn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L2PHIAn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L2PHIAn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L2PHIAn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIAn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIAn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L2PHIAn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIAn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIAn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L2PHIBn2_start                   : std_logic;
  signal VMSME_L2PHIBn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L2PHIBn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIBn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L2PHIBn2_wea          : t_VMSME_16_1b;
  signal VMSME_L2PHIBn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIBn2_din         : t_VMSME_16_DATA;
  signal VMSME_L2PHIBn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L2PHIBn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L2PHIBn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L2PHIBn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L2PHIBn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L2PHIBn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L2PHIBn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L2PHIBn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L2PHIBn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L2PHIBn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIBn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIBn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L2PHIBn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIBn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIBn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L2PHICn2_start                   : std_logic;
  signal VMSME_L2PHICn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L2PHICn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L2PHICn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L2PHICn2_wea          : t_VMSME_16_1b;
  signal VMSME_L2PHICn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L2PHICn2_din         : t_VMSME_16_DATA;
  signal VMSME_L2PHICn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L2PHICn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L2PHICn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L2PHICn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L2PHICn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L2PHICn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L2PHICn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L2PHICn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L2PHICn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L2PHICn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHICn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHICn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L2PHICn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHICn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHICn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L2PHIDn2_start                   : std_logic;
  signal VMSME_L2PHIDn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L2PHIDn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIDn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L2PHIDn2_wea          : t_VMSME_16_1b;
  signal VMSME_L2PHIDn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L2PHIDn2_din         : t_VMSME_16_DATA;
  signal VMSME_L2PHIDn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L2PHIDn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L2PHIDn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L2PHIDn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L2PHIDn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L2PHIDn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L2PHIDn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L2PHIDn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L2PHIDn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L2PHIDn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIDn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIDn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L2PHIDn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L2PHIDn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L2PHIDn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L3PHIAn2_start                   : std_logic;
  signal VMSME_L3PHIAn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L3PHIAn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIAn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L3PHIAn2_wea          : t_VMSME_16_1b;
  signal VMSME_L3PHIAn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIAn2_din         : t_VMSME_16_DATA;
  signal VMSME_L3PHIAn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L3PHIAn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L3PHIAn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L3PHIAn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L3PHIAn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L3PHIAn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L3PHIAn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L3PHIAn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L3PHIAn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L3PHIAn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIAn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIAn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L3PHIAn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIAn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIAn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L3PHIBn2_start                   : std_logic;
  signal VMSME_L3PHIBn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L3PHIBn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIBn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L3PHIBn2_wea          : t_VMSME_16_1b;
  signal VMSME_L3PHIBn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIBn2_din         : t_VMSME_16_DATA;
  signal VMSME_L3PHIBn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L3PHIBn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L3PHIBn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L3PHIBn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L3PHIBn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L3PHIBn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L3PHIBn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L3PHIBn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L3PHIBn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L3PHIBn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIBn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIBn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L3PHIBn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIBn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIBn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L3PHICn2_start                   : std_logic;
  signal VMSME_L3PHICn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L3PHICn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L3PHICn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L3PHICn2_wea          : t_VMSME_16_1b;
  signal VMSME_L3PHICn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L3PHICn2_din         : t_VMSME_16_DATA;
  signal VMSME_L3PHICn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L3PHICn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L3PHICn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L3PHICn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L3PHICn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L3PHICn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L3PHICn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L3PHICn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L3PHICn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L3PHICn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHICn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHICn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L3PHICn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHICn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHICn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L3PHIDn2_start                   : std_logic;
  signal VMSME_L3PHIDn2_wea_delay          : t_VMSME_16_1b;
  signal VMSME_L3PHIDn2_writeaddr_delay   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIDn2_din_delay         : t_VMSME_16_DATA;
  signal VMSME_L3PHIDn2_wea          : t_VMSME_16_1b;
  signal VMSME_L3PHIDn2_writeaddr   : t_VMSME_16_ADDR;
  signal VMSME_L3PHIDn2_din         : t_VMSME_16_DATA;
  signal VMSME_L3PHIDn2_A_enb         : t_VMSME_16_A1b;
  signal VMSME_L3PHIDn2_AV_readaddr   : t_VMSME_16_AADDR;
  signal VMSME_L3PHIDn2_AV_dout       : t_VMSME_16_ADATA;
  signal VMSME_L3PHIDn2_AV_dout_mask : t_VMSME_16_MASK; -- (#page)(#bin)
  signal VMSME_L3PHIDn2_enb_nent         : t_VMSME_16_1b;
  signal VMSME_L3PHIDn2_V_addr_nent   : t_VMSME_16_NENTADDR;
  signal VMSME_L3PHIDn2_AV_dout_nent : t_VMSME_16_NENT; -- (#page)(#bin)
  signal VMSME_L3PHIDn2_V_datatmp : t_VMSME_16_DATA_4;
  signal VMSME_L3PHIDn2_V_masktmp : t_VMSME_16_MASK_2;
  signal VMSME_L3PHIDn2_V_addr_binmaskA   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIDn2_V_binmaskA   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIDn2_enb_binmaskA   : t_VMSME_16_1b;
  signal VMSME_L3PHIDn2_V_addr_binmaskB   : t_VMSME_16_ADDRBINMASK;
  signal VMSME_L3PHIDn2_V_binmaskB   : t_VMSME_16_BINMASK;
  signal VMSME_L3PHIDn2_enb_binmaskB   : t_VMSME_16_1b;
  signal VMSME_L4PHIAn2_start                   : std_logic;
  signal VMSME_L4PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L4PHIAn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L4PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_L4PHIAn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_L4PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L4PHIAn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L4PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L4PHIAn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L4PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L4PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L4PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L4PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L4PHIAn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L4PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIAn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L4PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIAn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L4PHIBn2_start                   : std_logic;
  signal VMSME_L4PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L4PHIBn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L4PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_L4PHIBn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_L4PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L4PHIBn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L4PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L4PHIBn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L4PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L4PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L4PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L4PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L4PHIBn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L4PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIBn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L4PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIBn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L4PHICn2_start                   : std_logic;
  signal VMSME_L4PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L4PHICn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L4PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L4PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_L4PHICn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L4PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_L4PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L4PHICn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L4PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L4PHICn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L4PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L4PHICn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L4PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L4PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L4PHICn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L4PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHICn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L4PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHICn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L4PHIDn2_start                   : std_logic;
  signal VMSME_L4PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L4PHIDn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L4PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_L4PHIDn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L4PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_L4PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L4PHIDn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L4PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L4PHIDn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L4PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L4PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L4PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L4PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L4PHIDn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L4PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIDn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L4PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L4PHIDn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L4PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L5PHIAn2_start                   : std_logic;
  signal VMSME_L5PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L5PHIAn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L5PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_L5PHIAn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_L5PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L5PHIAn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L5PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L5PHIAn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L5PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L5PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L5PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L5PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L5PHIAn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L5PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIAn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L5PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIAn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L5PHIBn2_start                   : std_logic;
  signal VMSME_L5PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L5PHIBn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L5PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_L5PHIBn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_L5PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L5PHIBn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L5PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L5PHIBn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L5PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L5PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L5PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L5PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L5PHIBn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L5PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIBn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L5PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIBn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L5PHICn2_start                   : std_logic;
  signal VMSME_L5PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L5PHICn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L5PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L5PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_L5PHICn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L5PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_L5PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L5PHICn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L5PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L5PHICn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L5PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L5PHICn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L5PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L5PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L5PHICn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L5PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHICn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L5PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHICn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L5PHIDn2_start                   : std_logic;
  signal VMSME_L5PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L5PHIDn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L5PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_L5PHIDn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L5PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_L5PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L5PHIDn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L5PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L5PHIDn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L5PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L5PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L5PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L5PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L5PHIDn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L5PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIDn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L5PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L5PHIDn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L5PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L6PHIAn2_start                   : std_logic;
  signal VMSME_L6PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L6PHIAn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L6PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_L6PHIAn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_L6PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L6PHIAn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L6PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L6PHIAn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L6PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L6PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L6PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L6PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L6PHIAn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L6PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIAn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L6PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIAn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L6PHIBn2_start                   : std_logic;
  signal VMSME_L6PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L6PHIBn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L6PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_L6PHIBn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_L6PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L6PHIBn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L6PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L6PHIBn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L6PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L6PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L6PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L6PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L6PHIBn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L6PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIBn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L6PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIBn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L6PHICn2_start                   : std_logic;
  signal VMSME_L6PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L6PHICn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L6PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L6PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_L6PHICn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L6PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_L6PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L6PHICn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L6PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L6PHICn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L6PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L6PHICn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L6PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L6PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L6PHICn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L6PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHICn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L6PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHICn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_L6PHIDn2_start                   : std_logic;
  signal VMSME_L6PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_L6PHIDn2_writeaddr_delay   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_L6PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_L6PHIDn2_writeaddr   : t_VMSME_17_ADDR;
  signal VMSME_L6PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_L6PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_L6PHIDn2_AV_readaddr   : t_VMSME_17_AADDR;
  signal VMSME_L6PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_L6PHIDn2_AV_dout_mask : t_VMSME_17_MASK; -- (#page)(#bin)
  signal VMSME_L6PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_L6PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDR;
  signal VMSME_L6PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_L6PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_L6PHIDn2_V_masktmp : t_VMSME_17_MASK_2;
  signal VMSME_L6PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIDn2_V_binmaskA   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_L6PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASK;
  signal VMSME_L6PHIDn2_V_binmaskB   : t_VMSME_17_BINMASK;
  signal VMSME_L6PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D1PHIAn2_start                   : std_logic;
  signal VMSME_D1PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D1PHIAn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D1PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_D1PHIAn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_D1PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D1PHIAn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D1PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D1PHIAn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D1PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D1PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D1PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D1PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D1PHIAn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D1PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIAn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D1PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIAn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D1PHIBn2_start                   : std_logic;
  signal VMSME_D1PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D1PHIBn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D1PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_D1PHIBn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_D1PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D1PHIBn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D1PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D1PHIBn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D1PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D1PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D1PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D1PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D1PHIBn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D1PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIBn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D1PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIBn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D1PHICn2_start                   : std_logic;
  signal VMSME_D1PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D1PHICn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D1PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_D1PHICn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_D1PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D1PHICn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D1PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D1PHICn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D1PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D1PHICn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D1PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D1PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D1PHICn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D1PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHICn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D1PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHICn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D1PHIDn2_start                   : std_logic;
  signal VMSME_D1PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D1PHIDn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D1PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_D1PHIDn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D1PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_D1PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D1PHIDn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D1PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D1PHIDn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D1PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D1PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D1PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D1PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D1PHIDn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D1PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIDn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D1PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D1PHIDn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D1PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D2PHIAn2_start                   : std_logic;
  signal VMSME_D2PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D2PHIAn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D2PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_D2PHIAn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_D2PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D2PHIAn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D2PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D2PHIAn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D2PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D2PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D2PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D2PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D2PHIAn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D2PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIAn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D2PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIAn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D2PHIBn2_start                   : std_logic;
  signal VMSME_D2PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D2PHIBn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D2PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_D2PHIBn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_D2PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D2PHIBn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D2PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D2PHIBn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D2PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D2PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D2PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D2PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D2PHIBn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D2PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIBn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D2PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIBn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D2PHICn2_start                   : std_logic;
  signal VMSME_D2PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D2PHICn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D2PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_D2PHICn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_D2PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D2PHICn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D2PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D2PHICn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D2PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D2PHICn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D2PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D2PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D2PHICn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D2PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHICn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D2PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHICn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D2PHIDn2_start                   : std_logic;
  signal VMSME_D2PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D2PHIDn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D2PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_D2PHIDn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D2PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_D2PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D2PHIDn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D2PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D2PHIDn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D2PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D2PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D2PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D2PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D2PHIDn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D2PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIDn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D2PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D2PHIDn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D2PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D3PHIAn2_start                   : std_logic;
  signal VMSME_D3PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D3PHIAn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D3PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_D3PHIAn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_D3PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D3PHIAn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D3PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D3PHIAn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D3PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D3PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D3PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D3PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D3PHIAn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D3PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIAn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D3PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIAn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D3PHIBn2_start                   : std_logic;
  signal VMSME_D3PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D3PHIBn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D3PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_D3PHIBn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_D3PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D3PHIBn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D3PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D3PHIBn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D3PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D3PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D3PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D3PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D3PHIBn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D3PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIBn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D3PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIBn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D3PHICn2_start                   : std_logic;
  signal VMSME_D3PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D3PHICn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D3PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_D3PHICn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_D3PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D3PHICn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D3PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D3PHICn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D3PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D3PHICn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D3PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D3PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D3PHICn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D3PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHICn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D3PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHICn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D3PHIDn2_start                   : std_logic;
  signal VMSME_D3PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D3PHIDn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D3PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_D3PHIDn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D3PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_D3PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D3PHIDn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D3PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D3PHIDn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D3PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D3PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D3PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D3PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D3PHIDn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D3PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIDn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D3PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D3PHIDn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D3PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D4PHIAn2_start                   : std_logic;
  signal VMSME_D4PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D4PHIAn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D4PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_D4PHIAn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_D4PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D4PHIAn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D4PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D4PHIAn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D4PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D4PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D4PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D4PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D4PHIAn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D4PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIAn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D4PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIAn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D4PHIBn2_start                   : std_logic;
  signal VMSME_D4PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D4PHIBn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D4PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_D4PHIBn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_D4PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D4PHIBn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D4PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D4PHIBn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D4PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D4PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D4PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D4PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D4PHIBn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D4PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIBn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D4PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIBn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D4PHICn2_start                   : std_logic;
  signal VMSME_D4PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D4PHICn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D4PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_D4PHICn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_D4PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D4PHICn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D4PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D4PHICn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D4PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D4PHICn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D4PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D4PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D4PHICn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D4PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHICn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D4PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHICn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D4PHIDn2_start                   : std_logic;
  signal VMSME_D4PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D4PHIDn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D4PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_D4PHIDn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D4PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_D4PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D4PHIDn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D4PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D4PHIDn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D4PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D4PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D4PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D4PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D4PHIDn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D4PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIDn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D4PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D4PHIDn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D4PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D5PHIAn2_start                   : std_logic;
  signal VMSME_D5PHIAn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D5PHIAn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIAn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D5PHIAn2_wea          : t_VMSME_17_1b;
  signal VMSME_D5PHIAn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIAn2_din         : t_VMSME_17_DATA;
  signal VMSME_D5PHIAn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D5PHIAn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D5PHIAn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D5PHIAn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D5PHIAn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D5PHIAn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D5PHIAn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D5PHIAn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D5PHIAn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D5PHIAn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIAn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIAn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D5PHIAn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIAn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIAn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D5PHIBn2_start                   : std_logic;
  signal VMSME_D5PHIBn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D5PHIBn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIBn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D5PHIBn2_wea          : t_VMSME_17_1b;
  signal VMSME_D5PHIBn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIBn2_din         : t_VMSME_17_DATA;
  signal VMSME_D5PHIBn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D5PHIBn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D5PHIBn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D5PHIBn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D5PHIBn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D5PHIBn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D5PHIBn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D5PHIBn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D5PHIBn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D5PHIBn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIBn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIBn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D5PHIBn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIBn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIBn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D5PHICn2_start                   : std_logic;
  signal VMSME_D5PHICn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D5PHICn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHICn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D5PHICn2_wea          : t_VMSME_17_1b;
  signal VMSME_D5PHICn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHICn2_din         : t_VMSME_17_DATA;
  signal VMSME_D5PHICn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D5PHICn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D5PHICn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D5PHICn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D5PHICn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D5PHICn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D5PHICn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D5PHICn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D5PHICn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D5PHICn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHICn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHICn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D5PHICn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHICn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHICn2_enb_binmaskB   : t_VMSME_17_1b;
  signal VMSME_D5PHIDn2_start                   : std_logic;
  signal VMSME_D5PHIDn2_wea_delay          : t_VMSME_17_1b;
  signal VMSME_D5PHIDn2_writeaddr_delay   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIDn2_din_delay         : t_VMSME_17_DATA;
  signal VMSME_D5PHIDn2_wea          : t_VMSME_17_1b;
  signal VMSME_D5PHIDn2_writeaddr   : t_VMSME_17_ADDRDISK;
  signal VMSME_D5PHIDn2_din         : t_VMSME_17_DATA;
  signal VMSME_D5PHIDn2_A_enb         : t_VMSME_17_A1b;
  signal VMSME_D5PHIDn2_AV_readaddr   : t_VMSME_17_AADDRDISK;
  signal VMSME_D5PHIDn2_AV_dout       : t_VMSME_17_ADATA;
  signal VMSME_D5PHIDn2_AV_dout_mask : t_VMSME_17_MASKDISK; -- (#page)(#bin)
  signal VMSME_D5PHIDn2_enb_nent         : t_VMSME_17_1b;
  signal VMSME_D5PHIDn2_V_addr_nent   : t_VMSME_17_NENTADDRDISK;
  signal VMSME_D5PHIDn2_AV_dout_nent : t_VMSME_17_NENT; -- (#page)(#bin)
  signal VMSME_D5PHIDn2_V_datatmp : t_VMSME_17_DATA_4;
  signal VMSME_D5PHIDn2_V_masktmp : t_VMSME_17_MASKDISK_2;
  signal VMSME_D5PHIDn2_V_addr_binmaskA   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIDn2_V_binmaskA   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIDn2_enb_binmaskA   : t_VMSME_17_1b;
  signal VMSME_D5PHIDn2_V_addr_binmaskB   : t_VMSME_17_ADDRBINMASKDISK;
  signal VMSME_D5PHIDn2_V_binmaskB   : t_VMSME_17_BINMASKDISK;
  signal VMSME_D5PHIDn2_enb_binmaskB   : t_VMSME_17_1b;
  signal MPAR_L1L2ABCin_start                   : std_logic;
  signal MPAR_L1L2ABCin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2ABCin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2ABCin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2ABCin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2ABCin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2ABCin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2ABCin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2ABCin_valid        : STD_LOGIC;
  signal MPAR_L1L2ABCin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2ABCin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2ABCin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2DEin_start                   : std_logic;
  signal MPAR_L1L2DEin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2DEin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2DEin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2DEin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2DEin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2DEin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2DEin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2DEin_valid        : STD_LOGIC;
  signal MPAR_L1L2DEin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2DEin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2DEin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2Fin_start                   : std_logic;
  signal MPAR_L1L2Fin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2Fin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2Fin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2Fin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2Fin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2Fin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2Fin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2Fin_valid        : STD_LOGIC;
  signal MPAR_L1L2Fin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2Fin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2Fin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2Gin_start                   : std_logic;
  signal MPAR_L1L2Gin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2Gin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2Gin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2Gin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2Gin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2Gin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2Gin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2Gin_valid        : STD_LOGIC;
  signal MPAR_L1L2Gin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2Gin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2Gin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2HIin_start                   : std_logic;
  signal MPAR_L1L2HIin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2HIin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2HIin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2HIin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2HIin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2HIin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2HIin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2HIin_valid        : STD_LOGIC;
  signal MPAR_L1L2HIin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2HIin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2HIin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2JKLin_start                   : std_logic;
  signal MPAR_L1L2JKLin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2JKLin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2JKLin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2JKLin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2JKLin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2JKLin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2JKLin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1L2JKLin_valid        : STD_LOGIC;
  signal MPAR_L1L2JKLin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1L2JKLin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1L2JKLin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L2L3ABCDin_start                   : std_logic;
  signal MPAR_L2L3ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L2L3ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L2L3ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L2L3ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L2L3ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCDin_valid        : STD_LOGIC;
  signal MPAR_L2L3ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L2L3ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L2L3ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L3L4ABin_start                   : std_logic;
  signal MPAR_L3L4ABin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L3L4ABin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L3L4ABin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L3L4ABin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L3L4ABin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L3L4ABin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L3L4ABin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L3L4ABin_valid        : STD_LOGIC;
  signal MPAR_L3L4ABin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L3L4ABin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L3L4ABin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L3L4CDin_start                   : std_logic;
  signal MPAR_L3L4CDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L3L4CDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L3L4CDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L3L4CDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L3L4CDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L3L4CDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L3L4CDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L3L4CDin_valid        : STD_LOGIC;
  signal MPAR_L3L4CDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L3L4CDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L3L4CDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L5L6ABCDin_start                   : std_logic;
  signal MPAR_L5L6ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L5L6ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L5L6ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L5L6ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L5L6ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCDin_valid        : STD_LOGIC;
  signal MPAR_L5L6ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L5L6ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L5L6ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_D1D2ABCDin_start                   : std_logic;
  signal MPAR_D1D2ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_D1D2ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_D1D2ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_D1D2ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_D1D2ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCDin_valid        : STD_LOGIC;
  signal MPAR_D1D2ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_D1D2ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_D1D2ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_D3D4ABCDin_start                   : std_logic;
  signal MPAR_D3D4ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_D3D4ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_D3D4ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_D3D4ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_D3D4ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCDin_valid        : STD_LOGIC;
  signal MPAR_D3D4ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_D3D4ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_D3D4ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1D1ABCDin_start                   : std_logic;
  signal MPAR_L1D1ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1D1ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1D1ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1D1ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1D1ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCDin_valid        : STD_LOGIC;
  signal MPAR_L1D1ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1D1ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1D1ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1D1EFGHin_start                   : std_logic;
  signal MPAR_L1D1EFGHin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1D1EFGHin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1D1EFGHin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGHin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1D1EFGHin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1D1EFGHin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGHin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGHin_valid        : STD_LOGIC;
  signal MPAR_L1D1EFGHin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L1D1EFGHin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L1D1EFGHin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L2D1ABCDin_start                   : std_logic;
  signal MPAR_L2D1ABCDin_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L2D1ABCDin_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L2D1ABCDin_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCDin_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L2D1ABCDin_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L2D1ABCDin_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCDin_V_tpar        : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCDin_valid        : STD_LOGIC;
  signal MPAR_L2D1ABCDin_trackletindex        : STD_LOGIC_VECTOR(8 downto 0);
  signal MPAR_L2D1ABCDin_AV_dout_nent        : t_arr_7b(0 to 31);
  signal MPAR_L2D1ABCDin_AV_dout_mask        : t_arr_4b(0 to 7);
  signal MPAR_L1L2ABC_start                   : std_logic;
  signal MPAR_L1L2ABC_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2ABC_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2ABC_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2ABC_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2ABC_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2ABC_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2ABC_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2ABC_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2ABC_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2DE_start                   : std_logic;
  signal MPAR_L1L2DE_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2DE_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2DE_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2DE_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2DE_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2DE_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2DE_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2DE_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2DE_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2F_start                   : std_logic;
  signal MPAR_L1L2F_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2F_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2F_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2F_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2F_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2F_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2F_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2F_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2F_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2G_start                   : std_logic;
  signal MPAR_L1L2G_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2G_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2G_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2G_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2G_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2G_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2G_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2G_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2G_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2HI_start                   : std_logic;
  signal MPAR_L1L2HI_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2HI_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2HI_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2HI_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2HI_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2HI_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2HI_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2HI_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2HI_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1L2JKL_start                   : std_logic;
  signal MPAR_L1L2JKL_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1L2JKL_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1L2JKL_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1L2JKL_wea          : t_MPAR_73_1b;
  signal MPAR_L1L2JKL_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1L2JKL_din         : t_MPAR_73_DATA;
  signal MPAR_L1L2JKL_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1L2JKL_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1L2JKL_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCD_start                   : std_logic;
  signal MPAR_L2L3ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L2L3ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L2L3ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_L2L3ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L2L3ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_L2L3ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L2L3ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L2L3ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L3L4AB_start                   : std_logic;
  signal MPAR_L3L4AB_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L3L4AB_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L3L4AB_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L3L4AB_wea          : t_MPAR_73_1b;
  signal MPAR_L3L4AB_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L3L4AB_din         : t_MPAR_73_DATA;
  signal MPAR_L3L4AB_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L3L4AB_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L3L4AB_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L3L4CD_start                   : std_logic;
  signal MPAR_L3L4CD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L3L4CD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L3L4CD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L3L4CD_wea          : t_MPAR_73_1b;
  signal MPAR_L3L4CD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L3L4CD_din         : t_MPAR_73_DATA;
  signal MPAR_L3L4CD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L3L4CD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L3L4CD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCD_start                   : std_logic;
  signal MPAR_L5L6ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L5L6ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L5L6ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_L5L6ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L5L6ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_L5L6ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L5L6ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L5L6ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCD_start                   : std_logic;
  signal MPAR_D1D2ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_D1D2ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_D1D2ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_D1D2ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_D1D2ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_D1D2ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_D1D2ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_D1D2ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCD_start                   : std_logic;
  signal MPAR_D3D4ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_D3D4ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_D3D4ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_D3D4ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_D3D4ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_D3D4ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_D3D4ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_D3D4ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCD_start                   : std_logic;
  signal MPAR_L1D1ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1D1ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1D1ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_L1D1ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1D1ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_L1D1ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1D1ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1D1ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGH_start                   : std_logic;
  signal MPAR_L1D1EFGH_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L1D1EFGH_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L1D1EFGH_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGH_wea          : t_MPAR_73_1b;
  signal MPAR_L1D1EFGH_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L1D1EFGH_din         : t_MPAR_73_DATA;
  signal MPAR_L1D1EFGH_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L1D1EFGH_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L1D1EFGH_V_dout        : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCD_start                   : std_logic;
  signal MPAR_L2D1ABCD_wea_delay          : t_MPAR_73_1b;
  signal MPAR_L2D1ABCD_writeaddr_delay   : t_MPAR_73_ADDR;
  signal MPAR_L2D1ABCD_din_delay         : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCD_wea          : t_MPAR_73_1b;
  signal MPAR_L2D1ABCD_writeaddr   : t_MPAR_73_ADDR;
  signal MPAR_L2D1ABCD_din         : t_MPAR_73_DATA;
  signal MPAR_L2D1ABCD_enb          : t_MPAR_73_1b := '1';
  signal MPAR_L2D1ABCD_V_readaddr    : t_MPAR_73_ADDR;
  signal MPAR_L2D1ABCD_V_dout        : t_MPAR_73_DATA;
  signal MPROJ_L2L3ABCD_L1PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIA_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIA_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIA_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIA_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIB_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIB_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIB_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIB_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIC_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIC_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIC_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIC_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHID_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L1PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHID_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHID_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHID_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHID_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIE_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHIE_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L1PHIE_start                   : std_logic;
  signal MPROJ_L3L4CD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIE_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIE_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIE_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIE_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIE_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIE_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIE_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIE_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIE_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIE_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIE_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIE_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIE_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIE_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIF_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L1PHIF_start                   : std_logic;
  signal MPROJ_L3L4AB_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L1PHIF_start                   : std_logic;
  signal MPROJ_L3L4CD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIF_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIF_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIF_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIF_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIF_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIF_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIF_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIF_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIF_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIF_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIF_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIF_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIF_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIF_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIG_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L1PHIG_start                   : std_logic;
  signal MPROJ_L3L4CD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIG_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIG_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIG_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIG_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIG_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIG_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIG_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIG_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIG_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIG_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIG_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIG_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIG_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIG_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2L3ABCD_L1PHIH_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2L3ABCD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2L3ABCD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2L3ABCD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L1PHIH_start                   : std_logic;
  signal MPROJ_L3L4CD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L1PHIH_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L1PHIH_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D3D4ABCD_L1PHIH_start                   : std_logic;
  signal MPROJ_D3D4ABCD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_D3D4ABCD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D3D4ABCD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D3D4ABCD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L2D1ABCD_L1PHIH_start                   : std_logic;
  signal MPROJ_L2D1ABCD_L1PHIH_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIH_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIH_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIH_wea          : t_MPROJ_60_1b;
  signal MPROJ_L2D1ABCD_L1PHIH_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIH_din         : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIH_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L2D1ABCD_L1PHIH_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L2D1ABCD_L1PHIH_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_L1PHIH_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L2PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_L2PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L2PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L2PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L2PHIA_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L2PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L2PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L2PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L2PHIA_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L2PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L2PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L2PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L2PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_L2PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L2PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L2PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L2PHIB_start                   : std_logic;
  signal MPROJ_L3L4CD_L2PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L2PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L2PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L2PHIB_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L2PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L2PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L2PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L2PHIB_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L2PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L2PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L2PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4AB_L2PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_L2PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4AB_L2PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4AB_L2PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4AB_L2PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4AB_L2PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4AB_L2PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L2PHIC_start                   : std_logic;
  signal MPROJ_L3L4CD_L2PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L2PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L2PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L2PHIC_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L2PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L2PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L2PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L2PHIC_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L2PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L2PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L2PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L3L4CD_L2PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_L2PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L3L4CD_L2PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L3L4CD_L2PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L3L4CD_L2PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L3L4CD_L2PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L3L4CD_L2PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L2PHID_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L2PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L2PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L2PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L2PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L2PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L2PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_D1D2ABCD_L2PHID_start                   : std_logic;
  signal MPROJ_D1D2ABCD_L2PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_D1D2ABCD_L2PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_D1D2ABCD_L2PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_D1D2ABCD_L2PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_D1D2ABCD_L2PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_L2PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2ABC_L3PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_L3PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2ABC_L3PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2ABC_L3PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2ABC_L3PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L3PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2DE_L3PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_L3PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2DE_L3PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2DE_L3PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L3PHIA_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L3PHIA_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIA_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIA_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIA_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIA_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIA_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIA_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L3PHIA_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIA_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L3PHIA_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2ABC_L3PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2ABC_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2ABC_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2ABC_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2ABC_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2ABC_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2DE_L3PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2DE_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2DE_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2F_L3PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2F_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2F_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2F_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2F_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2G_L3PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2G_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2G_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2G_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2G_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2HI_L3PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2HI_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2HI_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L3PHIB_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L3PHIB_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIB_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIB_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIB_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIB_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIB_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIB_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L3PHIB_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIB_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L3PHIB_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2DE_L3PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2DE_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2DE_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2DE_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2DE_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2DE_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2F_L3PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2F_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2F_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2F_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2F_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2F_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2F_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2G_L3PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2G_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2G_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2G_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2G_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2G_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2G_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2HI_L3PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2HI_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2HI_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2JKL_L3PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2JKL_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2JKL_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2JKL_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L3PHIC_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L3PHIC_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIC_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIC_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIC_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHIC_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIC_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIC_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L3PHIC_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHIC_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L3PHIC_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2HI_L3PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_L3PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2HI_L3PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2HI_L3PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2HI_L3PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2HI_L3PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2HI_L3PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2JKL_L3PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_L3PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L1L2JKL_L3PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L1L2JKL_L3PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L1L2JKL_L3PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L1L2JKL_L3PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L1L2JKL_L3PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L3PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L5L6ABCD_L3PHID_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L3PHID_wea_delay          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHID_writeaddr_delay   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHID_din_delay         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHID_wea          : t_MPROJ_60_1b;
  signal MPROJ_L5L6ABCD_L3PHID_writeaddr   : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHID_din         : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHID_enb          : t_MPROJ_60_1b := '1';
  signal MPROJ_L5L6ABCD_L3PHID_V_readaddr    : t_MPROJ_60_ADDR;
  signal MPROJ_L5L6ABCD_L3PHID_V_dout        : t_MPROJ_60_DATA;
  signal MPROJ_L5L6ABCD_L3PHID_AV_dout_nent  : t_MPROJ_60_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L3PHID_AV_dout_mask  : t_MPROJ_60_MASK;
  signal MPROJ_L1L2ABC_L4PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_L4PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L4PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L4PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L4PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L4PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L4PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_L4PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L4PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L4PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L4PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_L4PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L4PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L4PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L4PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L4PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L4PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L4PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L5L6ABCD_L4PHIA_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L4PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L5L6ABCD_L4PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L4PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_L4PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L4PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L4PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L4PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L4PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L4PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L5L6ABCD_L4PHIB_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L4PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L5L6ABCD_L4PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L4PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L4PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L4PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L4PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L4PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L4PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L4PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L5L6ABCD_L4PHIC_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L4PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L5L6ABCD_L4PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L4PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L4PHID_start                   : std_logic;
  signal MPROJ_L1L2G_L4PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L4PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L4PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L4PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L4PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L4PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L4PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_L4PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L4PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L4PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L4PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L4PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L4PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L4PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_L4PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L4PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L4PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L4PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L4PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L4PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L4PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L4PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L4PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L4PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L4PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L4PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L4PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L4PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L5L6ABCD_L4PHID_start                   : std_logic;
  signal MPROJ_L5L6ABCD_L4PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L5L6ABCD_L4PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L5L6ABCD_L4PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L5L6ABCD_L4PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L5L6ABCD_L4PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L5L6ABCD_L4PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_L5PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_L5PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L5PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L5PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L5PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L5PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L5PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_L5PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L5PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L5PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L5PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_L5PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L5PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L5PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L5PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L5PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L5PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L5PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L5PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_L5PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L5PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L5PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_L5PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L5PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L5PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L5PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L5PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L5PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L5PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L5PHIB_start                   : std_logic;
  signal MPROJ_L3L4CD_L5PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L5PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L5PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L5PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L5PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L5PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L5PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L5PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L5PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L5PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L5PHIC_start                   : std_logic;
  signal MPROJ_L3L4CD_L5PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L5PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L5PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L5PHID_start                   : std_logic;
  signal MPROJ_L1L2G_L5PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L5PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L5PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L5PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L5PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L5PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L5PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_L5PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L5PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L5PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L5PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L5PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L5PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L5PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_L5PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L5PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L5PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L5PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L5PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L5PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L5PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L2L3ABCD_L5PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_L5PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L2L3ABCD_L5PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L2L3ABCD_L5PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L2L3ABCD_L5PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L2L3ABCD_L5PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_L5PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L5PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_L5PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L5PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L5PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L5PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L5PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L5PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_L6PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_L6PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L6PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L6PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L6PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L6PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L6PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_L6PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L6PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L6PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L6PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_L6PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L6PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L6PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L6PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_L6PHIA_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIA_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIA_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIA_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIA_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIA_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIA_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L6PHIA_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIA_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIA_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L6PHIA_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_L6PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2ABC_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2ABC_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2ABC_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2ABC_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2ABC_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L6PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L6PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L6PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L6PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L6PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L6PHIB_start                   : std_logic;
  signal MPROJ_L3L4CD_L6PHIB_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHIB_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIB_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIB_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHIB_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIB_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIB_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L6PHIB_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIB_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIB_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L6PHIB_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2DE_L6PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2DE_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2DE_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2DE_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2DE_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2DE_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2F_L6PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2F_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2F_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2F_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2F_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2F_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L6PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L6PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L6PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4AB_L6PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4AB_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4AB_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4AB_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4AB_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4AB_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L6PHIC_start                   : std_logic;
  signal MPROJ_L3L4CD_L6PHIC_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHIC_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIC_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIC_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHIC_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIC_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIC_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L6PHIC_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHIC_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHIC_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L6PHIC_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2G_L6PHID_start                   : std_logic;
  signal MPROJ_L1L2G_L6PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2G_L6PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2G_L6PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2G_L6PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2G_L6PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2G_L6PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2HI_L6PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_L6PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2HI_L6PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2HI_L6PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2HI_L6PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2HI_L6PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2HI_L6PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2JKL_L6PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_L6PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L6PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L1L2JKL_L6PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L1L2JKL_L6PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L1L2JKL_L6PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L1L2JKL_L6PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L1L2JKL_L6PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L3L4CD_L6PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_L6PHID_wea_delay          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHID_writeaddr_delay   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHID_din_delay         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHID_wea          : t_MPROJ_58_1b;
  signal MPROJ_L3L4CD_L6PHID_writeaddr   : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHID_din         : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHID_enb          : t_MPROJ_58_1b := '1';
  signal MPROJ_L3L4CD_L6PHID_V_readaddr    : t_MPROJ_58_ADDR;
  signal MPROJ_L3L4CD_L6PHID_V_dout        : t_MPROJ_58_DATA;
  signal MPROJ_L3L4CD_L6PHID_AV_dout_nent  : t_MPROJ_58_NENT; -- (#page)
  signal MPROJ_L3L4CD_L6PHID_AV_dout_mask  : t_MPROJ_58_MASK;
  signal MPROJ_L1L2ABC_D1PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D1PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D1PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D1PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D1PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D1PHIA_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D1PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D1PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D1PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D1PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D1PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D1PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D1PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D1PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D1PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D1PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D1PHIB_start                   : std_logic;
  signal MPROJ_L3L4CD_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D1PHIB_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D1PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D1PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D1PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D1PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D1PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D1PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D1PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D1PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D1PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D1PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D1PHIC_start                   : std_logic;
  signal MPROJ_L3L4CD_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D1PHIC_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D1PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D1PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D1PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D1PHID_start                   : std_logic;
  signal MPROJ_L1L2G_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D1PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D1PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D1PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D1PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D1PHID_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D1PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D1PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D1PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D1PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D1PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D1PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D2PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D2PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D2PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D2PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D2PHIA_start                   : std_logic;
  signal MPROJ_L3L4AB_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D2PHIA_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D2PHIA_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D2PHIA_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D2PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D2PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D2PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D2PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D2PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D2PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D2PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D2PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D2PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D2PHIB_start                   : std_logic;
  signal MPROJ_L3L4AB_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D2PHIB_start                   : std_logic;
  signal MPROJ_L3L4CD_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D2PHIB_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D2PHIB_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D2PHIB_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D2PHIB_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D2PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D2PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D2PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D2PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D2PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D2PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D2PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D2PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D2PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4AB_D2PHIC_start                   : std_logic;
  signal MPROJ_L3L4AB_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4AB_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4AB_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4AB_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4AB_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4AB_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D2PHIC_start                   : std_logic;
  signal MPROJ_L3L4CD_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D2PHIC_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D2PHIC_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D2PHIC_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D2PHIC_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D2PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D2PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D2PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D2PHID_start                   : std_logic;
  signal MPROJ_L1L2G_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D2PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D2PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D2PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L3L4CD_D2PHID_start                   : std_logic;
  signal MPROJ_L3L4CD_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L3L4CD_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L3L4CD_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L3L4CD_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L3L4CD_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L3L4CD_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D2PHID_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D2PHID_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D2PHID_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D2PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D2PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D2PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D2PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D2PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D2PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D3PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D3PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D3PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D3PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D3PHIA_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D3PHIA_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D3PHIA_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D3PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D3PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D3PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D3PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D3PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D3PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D3PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D3PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D3PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D3PHIB_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D3PHIB_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D3PHIB_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D3PHIB_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D3PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D3PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D3PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D3PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D3PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D3PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D3PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D3PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D3PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D3PHIC_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D3PHIC_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D3PHIC_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D3PHIC_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D3PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D3PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D3PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D3PHID_start                   : std_logic;
  signal MPROJ_L1L2G_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D3PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D3PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D3PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D3PHID_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D3PHID_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D3PHID_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D3PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D3PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D3PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D3PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D3PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D3PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D4PHIA_start                   : std_logic;
  signal MPROJ_L1L2ABC_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D4PHIA_start                   : std_logic;
  signal MPROJ_L1L2DE_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D4PHIA_start                   : std_logic;
  signal MPROJ_L1L2F_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D4PHIA_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D4PHIA_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D4PHIA_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D4PHIA_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D4PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D4PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D4PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2ABC_D4PHIB_start                   : std_logic;
  signal MPROJ_L1L2ABC_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2ABC_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2ABC_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2ABC_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2ABC_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2ABC_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D4PHIB_start                   : std_logic;
  signal MPROJ_L1L2DE_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D4PHIB_start                   : std_logic;
  signal MPROJ_L1L2F_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D4PHIB_start                   : std_logic;
  signal MPROJ_L1L2G_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D4PHIB_start                   : std_logic;
  signal MPROJ_L1L2HI_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D4PHIB_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D4PHIB_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D4PHIB_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D4PHIB_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D4PHIB_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D4PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D4PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D4PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2DE_D4PHIC_start                   : std_logic;
  signal MPROJ_L1L2DE_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2DE_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2DE_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2DE_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2DE_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2DE_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2F_D4PHIC_start                   : std_logic;
  signal MPROJ_L1L2F_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2F_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2F_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2F_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2F_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2F_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D4PHIC_start                   : std_logic;
  signal MPROJ_L1L2G_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D4PHIC_start                   : std_logic;
  signal MPROJ_L1L2HI_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D4PHIC_start                   : std_logic;
  signal MPROJ_L1L2JKL_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D4PHIC_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D4PHIC_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D4PHIC_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D4PHIC_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D4PHIC_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D4PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D4PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D4PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2G_D4PHID_start                   : std_logic;
  signal MPROJ_L1L2G_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2G_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2G_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2G_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2G_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2G_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2HI_D4PHID_start                   : std_logic;
  signal MPROJ_L1L2HI_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2HI_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2HI_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2HI_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2HI_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2HI_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1L2JKL_D4PHID_start                   : std_logic;
  signal MPROJ_L1L2JKL_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1L2JKL_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1L2JKL_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1L2JKL_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1L2JKL_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1L2JKL_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2L3ABCD_D4PHID_start                   : std_logic;
  signal MPROJ_L2L3ABCD_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2L3ABCD_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2L3ABCD_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2L3ABCD_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2L3ABCD_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2L3ABCD_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D4PHID_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D4PHID_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L2D1ABCD_D4PHID_start                   : std_logic;
  signal MPROJ_L2D1ABCD_D4PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L2D1ABCD_D4PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L2D1ABCD_D4PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L2D1ABCD_D4PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L2D1ABCD_D4PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L2D1ABCD_D4PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D5PHIA_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D5PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D5PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D5PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D5PHIA_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D5PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D5PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D5PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D5PHIA_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D5PHIA_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIA_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIA_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIA_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIA_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIA_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIA_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D5PHIA_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIA_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D5PHIA_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D5PHIB_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D5PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D5PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D5PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D5PHIB_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D5PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D5PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D5PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D5PHIB_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D5PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D5PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D5PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D5PHIB_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D5PHIB_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHIB_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIB_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIB_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHIB_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIB_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIB_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D5PHIB_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIB_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D5PHIB_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D5PHIC_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D5PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D5PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D5PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D5PHIC_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D5PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D5PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D5PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1ABCD_D5PHIC_start                   : std_logic;
  signal MPROJ_L1D1ABCD_D5PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1ABCD_D5PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1ABCD_D5PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1ABCD_D5PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1ABCD_D5PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D5PHIC_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D5PHIC_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHIC_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIC_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIC_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHIC_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIC_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIC_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D5PHIC_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHIC_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D5PHIC_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D1D2ABCD_D5PHID_start                   : std_logic;
  signal MPROJ_D1D2ABCD_D5PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D1D2ABCD_D5PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D1D2ABCD_D5PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D1D2ABCD_D5PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D1D2ABCD_D5PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D1D2ABCD_D5PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_D3D4ABCD_D5PHID_start                   : std_logic;
  signal MPROJ_D3D4ABCD_D5PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_D3D4ABCD_D5PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_D3D4ABCD_D5PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_D3D4ABCD_D5PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_D3D4ABCD_D5PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_D3D4ABCD_D5PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal MPROJ_L1D1EFGH_D5PHID_start                   : std_logic;
  signal MPROJ_L1D1EFGH_D5PHID_wea_delay          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHID_writeaddr_delay   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHID_din_delay         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHID_wea          : t_MPROJ_59_1b;
  signal MPROJ_L1D1EFGH_D5PHID_writeaddr   : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHID_din         : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHID_enb          : t_MPROJ_59_1b := '1';
  signal MPROJ_L1D1EFGH_D5PHID_V_readaddr    : t_MPROJ_59_ADDR;
  signal MPROJ_L1D1EFGH_D5PHID_V_dout        : t_MPROJ_59_DATA;
  signal MPROJ_L1D1EFGH_D5PHID_AV_dout_nent  : t_MPROJ_59_NENT; -- (#page)
  signal MPROJ_L1D1EFGH_D5PHID_AV_dout_mask  : t_MPROJ_59_MASK;
  signal FM_AAAA_L1PHIA_start                   : std_logic;
  signal FM_AAAA_L1PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIA_start                   : std_logic;
  signal FM_BBBB_L1PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIB_start                   : std_logic;
  signal FM_AAAA_L1PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIB_start                   : std_logic;
  signal FM_BBBB_L1PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIC_start                   : std_logic;
  signal FM_AAAA_L1PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIC_start                   : std_logic;
  signal FM_BBBB_L1PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHID_start                   : std_logic;
  signal FM_AAAA_L1PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHID_start                   : std_logic;
  signal FM_BBBB_L1PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIE_start                   : std_logic;
  signal FM_AAAA_L1PHIE_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIE_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIE_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIE_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIE_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIE_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIE_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIE_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIE_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIE_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIE_start                   : std_logic;
  signal FM_BBBB_L1PHIE_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIE_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIE_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIE_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIE_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIE_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIE_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIE_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIE_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIE_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIF_start                   : std_logic;
  signal FM_AAAA_L1PHIF_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIF_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIF_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIF_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIF_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIF_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIF_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIF_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIF_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIF_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIF_start                   : std_logic;
  signal FM_BBBB_L1PHIF_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIF_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIF_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIF_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIF_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIF_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIF_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIF_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIF_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIF_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIG_start                   : std_logic;
  signal FM_AAAA_L1PHIG_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIG_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIG_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIG_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIG_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIG_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIG_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIG_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIG_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIG_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIG_start                   : std_logic;
  signal FM_BBBB_L1PHIG_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIG_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIG_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIG_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIG_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIG_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIG_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIG_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIG_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIG_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L1PHIH_start                   : std_logic;
  signal FM_AAAA_L1PHIH_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L1PHIH_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIH_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIH_wea          : t_FM_52_1b;
  signal FM_AAAA_L1PHIH_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIH_din         : t_FM_52_DATA;
  signal FM_AAAA_L1PHIH_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L1PHIH_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L1PHIH_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L1PHIH_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L1PHIH_start                   : std_logic;
  signal FM_BBBB_L1PHIH_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L1PHIH_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIH_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIH_wea          : t_FM_52_1b;
  signal FM_BBBB_L1PHIH_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIH_din         : t_FM_52_DATA;
  signal FM_BBBB_L1PHIH_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L1PHIH_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L1PHIH_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L1PHIH_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L2PHIA_start                   : std_logic;
  signal FM_AAAA_L2PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L2PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L2PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L2PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L2PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L2PHIA_start                   : std_logic;
  signal FM_BBBB_L2PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L2PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L2PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L2PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L2PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L2PHIB_start                   : std_logic;
  signal FM_AAAA_L2PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L2PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L2PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L2PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L2PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L2PHIB_start                   : std_logic;
  signal FM_BBBB_L2PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L2PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L2PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L2PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L2PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L2PHIC_start                   : std_logic;
  signal FM_AAAA_L2PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L2PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L2PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L2PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L2PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L2PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L2PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L2PHIC_start                   : std_logic;
  signal FM_BBBB_L2PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L2PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L2PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L2PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L2PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L2PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L2PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L2PHID_start                   : std_logic;
  signal FM_AAAA_L2PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L2PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L2PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L2PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L2PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L2PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L2PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L2PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L2PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L2PHID_start                   : std_logic;
  signal FM_BBBB_L2PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L2PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L2PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L2PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L2PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L2PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L2PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L2PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L2PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L3PHIA_start                   : std_logic;
  signal FM_AAAA_L3PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L3PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L3PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L3PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L3PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L3PHIA_start                   : std_logic;
  signal FM_BBBB_L3PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L3PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L3PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L3PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L3PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L3PHIB_start                   : std_logic;
  signal FM_AAAA_L3PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L3PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L3PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L3PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L3PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L3PHIB_start                   : std_logic;
  signal FM_BBBB_L3PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L3PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L3PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L3PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L3PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L3PHIC_start                   : std_logic;
  signal FM_AAAA_L3PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L3PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L3PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L3PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L3PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L3PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L3PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L3PHIC_start                   : std_logic;
  signal FM_BBBB_L3PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L3PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L3PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L3PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L3PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L3PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L3PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L3PHID_start                   : std_logic;
  signal FM_AAAA_L3PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L3PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L3PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L3PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L3PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L3PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L3PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L3PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L3PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L3PHID_start                   : std_logic;
  signal FM_BBBB_L3PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L3PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L3PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L3PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L3PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L3PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L3PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L3PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L3PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L4PHIA_start                   : std_logic;
  signal FM_AAAA_L4PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L4PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L4PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L4PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L4PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L4PHIA_start                   : std_logic;
  signal FM_BBBB_L4PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L4PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L4PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L4PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L4PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L4PHIB_start                   : std_logic;
  signal FM_AAAA_L4PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L4PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L4PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L4PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L4PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L4PHIB_start                   : std_logic;
  signal FM_BBBB_L4PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L4PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L4PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L4PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L4PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L4PHIC_start                   : std_logic;
  signal FM_AAAA_L4PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L4PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L4PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L4PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L4PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L4PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L4PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L4PHIC_start                   : std_logic;
  signal FM_BBBB_L4PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L4PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L4PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L4PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L4PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L4PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L4PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L4PHID_start                   : std_logic;
  signal FM_AAAA_L4PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L4PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L4PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L4PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L4PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L4PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L4PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L4PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L4PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L4PHID_start                   : std_logic;
  signal FM_BBBB_L4PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L4PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L4PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L4PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L4PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L4PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L4PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L4PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L4PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L5PHIA_start                   : std_logic;
  signal FM_AAAA_L5PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L5PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L5PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L5PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L5PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L5PHIA_start                   : std_logic;
  signal FM_BBBB_L5PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L5PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L5PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L5PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L5PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L5PHIB_start                   : std_logic;
  signal FM_AAAA_L5PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L5PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L5PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L5PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L5PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L5PHIB_start                   : std_logic;
  signal FM_BBBB_L5PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L5PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L5PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L5PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L5PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L5PHIC_start                   : std_logic;
  signal FM_AAAA_L5PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L5PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L5PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L5PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L5PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L5PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L5PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L5PHIC_start                   : std_logic;
  signal FM_BBBB_L5PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L5PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L5PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L5PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L5PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L5PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L5PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L5PHID_start                   : std_logic;
  signal FM_AAAA_L5PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L5PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L5PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L5PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L5PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L5PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L5PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L5PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L5PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L5PHID_start                   : std_logic;
  signal FM_BBBB_L5PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L5PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L5PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L5PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L5PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L5PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L5PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L5PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L5PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L6PHIA_start                   : std_logic;
  signal FM_AAAA_L6PHIA_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L6PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIA_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIA_wea          : t_FM_52_1b;
  signal FM_AAAA_L6PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIA_din         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIA_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L6PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIA_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L6PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L6PHIA_start                   : std_logic;
  signal FM_BBBB_L6PHIA_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L6PHIA_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIA_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIA_wea          : t_FM_52_1b;
  signal FM_BBBB_L6PHIA_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIA_din         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIA_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L6PHIA_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIA_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L6PHIA_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L6PHIB_start                   : std_logic;
  signal FM_AAAA_L6PHIB_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L6PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIB_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIB_wea          : t_FM_52_1b;
  signal FM_AAAA_L6PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIB_din         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIB_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L6PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIB_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L6PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L6PHIB_start                   : std_logic;
  signal FM_BBBB_L6PHIB_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L6PHIB_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIB_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIB_wea          : t_FM_52_1b;
  signal FM_BBBB_L6PHIB_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIB_din         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIB_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L6PHIB_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIB_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L6PHIB_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L6PHIC_start                   : std_logic;
  signal FM_AAAA_L6PHIC_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L6PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIC_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIC_wea          : t_FM_52_1b;
  signal FM_AAAA_L6PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIC_din         : t_FM_52_DATA;
  signal FM_AAAA_L6PHIC_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L6PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L6PHIC_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L6PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L6PHIC_start                   : std_logic;
  signal FM_BBBB_L6PHIC_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L6PHIC_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIC_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIC_wea          : t_FM_52_1b;
  signal FM_BBBB_L6PHIC_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIC_din         : t_FM_52_DATA;
  signal FM_BBBB_L6PHIC_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L6PHIC_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L6PHIC_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L6PHIC_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_L6PHID_start                   : std_logic;
  signal FM_AAAA_L6PHID_wea_delay          : t_FM_52_1b;
  signal FM_AAAA_L6PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHID_din_delay         : t_FM_52_DATA;
  signal FM_AAAA_L6PHID_wea          : t_FM_52_1b;
  signal FM_AAAA_L6PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_AAAA_L6PHID_din         : t_FM_52_DATA;
  signal FM_AAAA_L6PHID_enb          : t_FM_52_1b := '1';
  signal FM_AAAA_L6PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_AAAA_L6PHID_V_dout        : t_FM_52_DATA;
  signal FM_AAAA_L6PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_BBBB_L6PHID_start                   : std_logic;
  signal FM_BBBB_L6PHID_wea_delay          : t_FM_52_1b;
  signal FM_BBBB_L6PHID_writeaddr_delay   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHID_din_delay         : t_FM_52_DATA;
  signal FM_BBBB_L6PHID_wea          : t_FM_52_1b;
  signal FM_BBBB_L6PHID_writeaddr   : t_FM_52_ADDR;
  signal FM_BBBB_L6PHID_din         : t_FM_52_DATA;
  signal FM_BBBB_L6PHID_enb          : t_FM_52_1b := '1';
  signal FM_BBBB_L6PHID_V_readaddr    : t_FM_52_ADDR;
  signal FM_BBBB_L6PHID_V_dout        : t_FM_52_DATA;
  signal FM_BBBB_L6PHID_AV_dout_nent  : t_FM_52_NENT; -- (#page)
  signal FM_AAAA_D1PHIA_start                   : std_logic;
  signal FM_AAAA_D1PHIA_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D1PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIA_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIA_wea          : t_FM_55_1b;
  signal FM_AAAA_D1PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIA_din         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIA_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D1PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIA_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D1PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D1PHIA_start                   : std_logic;
  signal FM_BBBB_D1PHIA_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D1PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIA_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIA_wea          : t_FM_55_1b;
  signal FM_BBBB_D1PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIA_din         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIA_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D1PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIA_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D1PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D1PHIB_start                   : std_logic;
  signal FM_AAAA_D1PHIB_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D1PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIB_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIB_wea          : t_FM_55_1b;
  signal FM_AAAA_D1PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIB_din         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIB_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D1PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIB_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D1PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D1PHIB_start                   : std_logic;
  signal FM_BBBB_D1PHIB_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D1PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIB_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIB_wea          : t_FM_55_1b;
  signal FM_BBBB_D1PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIB_din         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIB_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D1PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIB_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D1PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D1PHIC_start                   : std_logic;
  signal FM_AAAA_D1PHIC_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D1PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIC_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIC_wea          : t_FM_55_1b;
  signal FM_AAAA_D1PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIC_din         : t_FM_55_DATA;
  signal FM_AAAA_D1PHIC_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D1PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D1PHIC_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D1PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D1PHIC_start                   : std_logic;
  signal FM_BBBB_D1PHIC_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D1PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIC_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIC_wea          : t_FM_55_1b;
  signal FM_BBBB_D1PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIC_din         : t_FM_55_DATA;
  signal FM_BBBB_D1PHIC_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D1PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D1PHIC_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D1PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D1PHID_start                   : std_logic;
  signal FM_AAAA_D1PHID_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D1PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHID_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D1PHID_wea          : t_FM_55_1b;
  signal FM_AAAA_D1PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D1PHID_din         : t_FM_55_DATA;
  signal FM_AAAA_D1PHID_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D1PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D1PHID_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D1PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D1PHID_start                   : std_logic;
  signal FM_BBBB_D1PHID_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D1PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHID_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D1PHID_wea          : t_FM_55_1b;
  signal FM_BBBB_D1PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D1PHID_din         : t_FM_55_DATA;
  signal FM_BBBB_D1PHID_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D1PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D1PHID_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D1PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D2PHIA_start                   : std_logic;
  signal FM_AAAA_D2PHIA_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D2PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIA_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIA_wea          : t_FM_55_1b;
  signal FM_AAAA_D2PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIA_din         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIA_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D2PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIA_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D2PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D2PHIA_start                   : std_logic;
  signal FM_BBBB_D2PHIA_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D2PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIA_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIA_wea          : t_FM_55_1b;
  signal FM_BBBB_D2PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIA_din         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIA_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D2PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIA_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D2PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D2PHIB_start                   : std_logic;
  signal FM_AAAA_D2PHIB_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D2PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIB_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIB_wea          : t_FM_55_1b;
  signal FM_AAAA_D2PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIB_din         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIB_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D2PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIB_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D2PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D2PHIB_start                   : std_logic;
  signal FM_BBBB_D2PHIB_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D2PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIB_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIB_wea          : t_FM_55_1b;
  signal FM_BBBB_D2PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIB_din         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIB_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D2PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIB_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D2PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D2PHIC_start                   : std_logic;
  signal FM_AAAA_D2PHIC_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D2PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIC_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIC_wea          : t_FM_55_1b;
  signal FM_AAAA_D2PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIC_din         : t_FM_55_DATA;
  signal FM_AAAA_D2PHIC_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D2PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D2PHIC_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D2PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D2PHIC_start                   : std_logic;
  signal FM_BBBB_D2PHIC_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D2PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIC_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIC_wea          : t_FM_55_1b;
  signal FM_BBBB_D2PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIC_din         : t_FM_55_DATA;
  signal FM_BBBB_D2PHIC_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D2PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D2PHIC_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D2PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D2PHID_start                   : std_logic;
  signal FM_AAAA_D2PHID_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D2PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHID_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D2PHID_wea          : t_FM_55_1b;
  signal FM_AAAA_D2PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D2PHID_din         : t_FM_55_DATA;
  signal FM_AAAA_D2PHID_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D2PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D2PHID_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D2PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D2PHID_start                   : std_logic;
  signal FM_BBBB_D2PHID_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D2PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHID_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D2PHID_wea          : t_FM_55_1b;
  signal FM_BBBB_D2PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D2PHID_din         : t_FM_55_DATA;
  signal FM_BBBB_D2PHID_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D2PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D2PHID_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D2PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D3PHIA_start                   : std_logic;
  signal FM_AAAA_D3PHIA_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D3PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIA_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIA_wea          : t_FM_55_1b;
  signal FM_AAAA_D3PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIA_din         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIA_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D3PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIA_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D3PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D3PHIA_start                   : std_logic;
  signal FM_BBBB_D3PHIA_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D3PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIA_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIA_wea          : t_FM_55_1b;
  signal FM_BBBB_D3PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIA_din         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIA_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D3PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIA_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D3PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D3PHIB_start                   : std_logic;
  signal FM_AAAA_D3PHIB_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D3PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIB_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIB_wea          : t_FM_55_1b;
  signal FM_AAAA_D3PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIB_din         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIB_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D3PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIB_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D3PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D3PHIB_start                   : std_logic;
  signal FM_BBBB_D3PHIB_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D3PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIB_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIB_wea          : t_FM_55_1b;
  signal FM_BBBB_D3PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIB_din         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIB_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D3PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIB_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D3PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D3PHIC_start                   : std_logic;
  signal FM_AAAA_D3PHIC_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D3PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIC_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIC_wea          : t_FM_55_1b;
  signal FM_AAAA_D3PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIC_din         : t_FM_55_DATA;
  signal FM_AAAA_D3PHIC_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D3PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D3PHIC_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D3PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D3PHIC_start                   : std_logic;
  signal FM_BBBB_D3PHIC_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D3PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIC_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIC_wea          : t_FM_55_1b;
  signal FM_BBBB_D3PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIC_din         : t_FM_55_DATA;
  signal FM_BBBB_D3PHIC_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D3PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D3PHIC_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D3PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D3PHID_start                   : std_logic;
  signal FM_AAAA_D3PHID_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D3PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHID_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D3PHID_wea          : t_FM_55_1b;
  signal FM_AAAA_D3PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D3PHID_din         : t_FM_55_DATA;
  signal FM_AAAA_D3PHID_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D3PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D3PHID_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D3PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D3PHID_start                   : std_logic;
  signal FM_BBBB_D3PHID_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D3PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHID_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D3PHID_wea          : t_FM_55_1b;
  signal FM_BBBB_D3PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D3PHID_din         : t_FM_55_DATA;
  signal FM_BBBB_D3PHID_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D3PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D3PHID_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D3PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D4PHIA_start                   : std_logic;
  signal FM_AAAA_D4PHIA_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D4PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIA_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIA_wea          : t_FM_55_1b;
  signal FM_AAAA_D4PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIA_din         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIA_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D4PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIA_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D4PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D4PHIA_start                   : std_logic;
  signal FM_BBBB_D4PHIA_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D4PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIA_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIA_wea          : t_FM_55_1b;
  signal FM_BBBB_D4PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIA_din         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIA_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D4PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIA_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D4PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D4PHIB_start                   : std_logic;
  signal FM_AAAA_D4PHIB_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D4PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIB_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIB_wea          : t_FM_55_1b;
  signal FM_AAAA_D4PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIB_din         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIB_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D4PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIB_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D4PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D4PHIB_start                   : std_logic;
  signal FM_BBBB_D4PHIB_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D4PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIB_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIB_wea          : t_FM_55_1b;
  signal FM_BBBB_D4PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIB_din         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIB_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D4PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIB_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D4PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D4PHIC_start                   : std_logic;
  signal FM_AAAA_D4PHIC_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D4PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIC_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIC_wea          : t_FM_55_1b;
  signal FM_AAAA_D4PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIC_din         : t_FM_55_DATA;
  signal FM_AAAA_D4PHIC_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D4PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D4PHIC_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D4PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D4PHIC_start                   : std_logic;
  signal FM_BBBB_D4PHIC_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D4PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIC_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIC_wea          : t_FM_55_1b;
  signal FM_BBBB_D4PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIC_din         : t_FM_55_DATA;
  signal FM_BBBB_D4PHIC_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D4PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D4PHIC_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D4PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D4PHID_start                   : std_logic;
  signal FM_AAAA_D4PHID_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D4PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHID_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D4PHID_wea          : t_FM_55_1b;
  signal FM_AAAA_D4PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D4PHID_din         : t_FM_55_DATA;
  signal FM_AAAA_D4PHID_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D4PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D4PHID_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D4PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D4PHID_start                   : std_logic;
  signal FM_BBBB_D4PHID_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D4PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHID_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D4PHID_wea          : t_FM_55_1b;
  signal FM_BBBB_D4PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D4PHID_din         : t_FM_55_DATA;
  signal FM_BBBB_D4PHID_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D4PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D4PHID_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D4PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D5PHIA_start                   : std_logic;
  signal FM_AAAA_D5PHIA_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D5PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIA_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIA_wea          : t_FM_55_1b;
  signal FM_AAAA_D5PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIA_din         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIA_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D5PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIA_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D5PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D5PHIA_start                   : std_logic;
  signal FM_BBBB_D5PHIA_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D5PHIA_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIA_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIA_wea          : t_FM_55_1b;
  signal FM_BBBB_D5PHIA_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIA_din         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIA_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D5PHIA_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIA_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D5PHIA_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D5PHIB_start                   : std_logic;
  signal FM_AAAA_D5PHIB_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D5PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIB_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIB_wea          : t_FM_55_1b;
  signal FM_AAAA_D5PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIB_din         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIB_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D5PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIB_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D5PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D5PHIB_start                   : std_logic;
  signal FM_BBBB_D5PHIB_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D5PHIB_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIB_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIB_wea          : t_FM_55_1b;
  signal FM_BBBB_D5PHIB_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIB_din         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIB_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D5PHIB_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIB_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D5PHIB_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D5PHIC_start                   : std_logic;
  signal FM_AAAA_D5PHIC_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D5PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIC_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIC_wea          : t_FM_55_1b;
  signal FM_AAAA_D5PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIC_din         : t_FM_55_DATA;
  signal FM_AAAA_D5PHIC_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D5PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D5PHIC_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D5PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D5PHIC_start                   : std_logic;
  signal FM_BBBB_D5PHIC_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D5PHIC_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIC_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIC_wea          : t_FM_55_1b;
  signal FM_BBBB_D5PHIC_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIC_din         : t_FM_55_DATA;
  signal FM_BBBB_D5PHIC_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D5PHIC_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D5PHIC_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D5PHIC_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_AAAA_D5PHID_start                   : std_logic;
  signal FM_AAAA_D5PHID_wea_delay          : t_FM_55_1b;
  signal FM_AAAA_D5PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHID_din_delay         : t_FM_55_DATA;
  signal FM_AAAA_D5PHID_wea          : t_FM_55_1b;
  signal FM_AAAA_D5PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_AAAA_D5PHID_din         : t_FM_55_DATA;
  signal FM_AAAA_D5PHID_enb          : t_FM_55_1b := '1';
  signal FM_AAAA_D5PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_AAAA_D5PHID_V_dout        : t_FM_55_DATA;
  signal FM_AAAA_D5PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal FM_BBBB_D5PHID_start                   : std_logic;
  signal FM_BBBB_D5PHID_wea_delay          : t_FM_55_1b;
  signal FM_BBBB_D5PHID_writeaddr_delay   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHID_din_delay         : t_FM_55_DATA;
  signal FM_BBBB_D5PHID_wea          : t_FM_55_1b;
  signal FM_BBBB_D5PHID_writeaddr   : t_FM_55_ADDR;
  signal FM_BBBB_D5PHID_din         : t_FM_55_DATA;
  signal FM_BBBB_D5PHID_enb          : t_FM_55_1b := '1';
  signal FM_BBBB_D5PHID_V_readaddr    : t_FM_55_ADDR;
  signal FM_BBBB_D5PHID_V_dout        : t_FM_55_DATA;
  signal FM_BBBB_D5PHID_AV_dout_nent  : t_FM_55_NENT; -- (#page)
  signal VMSMER_L1PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIA_start : std_logic := '0';
  signal VMSMER_L1PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIB_start : std_logic := '0';
  signal VMSMER_L1PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIC_start : std_logic := '0';
  signal VMSMER_L1PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHID_start : std_logic := '0';
  signal VMSMER_L1PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIE_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIE_start : std_logic := '0';
  signal VMSMER_L1PHIE_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIF_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIF_start : std_logic := '0';
  signal VMSMER_L1PHIF_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIG_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIG_start : std_logic := '0';
  signal VMSMER_L1PHIG_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIH_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L1PHIH_start : std_logic := '0';
  signal VMSMER_L1PHIH_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIA_start : std_logic := '0';
  signal VMSMER_L2PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIB_start : std_logic := '0';
  signal VMSMER_L2PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHIC_start : std_logic := '0';
  signal VMSMER_L2PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L2PHID_start : std_logic := '0';
  signal VMSMER_L2PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIA_start : std_logic := '0';
  signal VMSMER_L3PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIB_start : std_logic := '0';
  signal VMSMER_L3PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHIC_start : std_logic := '0';
  signal VMSMER_L3PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L3PHID_start : std_logic := '0';
  signal VMSMER_L3PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIA_start : std_logic := '0';
  signal VMSMER_L4PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIB_start : std_logic := '0';
  signal VMSMER_L4PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHIC_start : std_logic := '0';
  signal VMSMER_L4PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L4PHID_start : std_logic := '0';
  signal VMSMER_L4PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIA_start : std_logic := '0';
  signal VMSMER_L5PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIB_start : std_logic := '0';
  signal VMSMER_L5PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHIC_start : std_logic := '0';
  signal VMSMER_L5PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L5PHID_start : std_logic := '0';
  signal VMSMER_L5PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIA_start : std_logic := '0';
  signal VMSMER_L6PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIB_start : std_logic := '0';
  signal VMSMER_L6PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHIC_start : std_logic := '0';
  signal VMSMER_L6PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_L6PHID_start : std_logic := '0';
  signal VMSMER_L6PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIA_start : std_logic := '0';
  signal VMSMER_D1PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIB_start : std_logic := '0';
  signal VMSMER_D1PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHIC_start : std_logic := '0';
  signal VMSMER_D1PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D1PHID_start : std_logic := '0';
  signal VMSMER_D1PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIA_start : std_logic := '0';
  signal VMSMER_D2PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIB_start : std_logic := '0';
  signal VMSMER_D2PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHIC_start : std_logic := '0';
  signal VMSMER_D2PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D2PHID_start : std_logic := '0';
  signal VMSMER_D2PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIA_start : std_logic := '0';
  signal VMSMER_D3PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIB_start : std_logic := '0';
  signal VMSMER_D3PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHIC_start : std_logic := '0';
  signal VMSMER_D3PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D3PHID_start : std_logic := '0';
  signal VMSMER_D3PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIA_start : std_logic := '0';
  signal VMSMER_D4PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIB_start : std_logic := '0';
  signal VMSMER_D4PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHIC_start : std_logic := '0';
  signal VMSMER_D4PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D4PHID_start : std_logic := '0';
  signal VMSMER_D4PHID_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIA_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIA_start : std_logic := '0';
  signal VMSMER_D5PHIA_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIB_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIB_start : std_logic := '0';
  signal VMSMER_D5PHIB_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIC_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHIC_start : std_logic := '0';
  signal VMSMER_D5PHIC_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHID_bx : std_logic_vector(2 downto 0);
  signal VMSMER_D5PHID_start : std_logic := '0';
  signal VMSMER_D5PHID_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2ABC_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2ABC_start : std_logic := '0';
  signal PC_L1L2ABC_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2DE_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2DE_start : std_logic := '0';
  signal PC_L1L2DE_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2F_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2F_start : std_logic := '0';
  signal PC_L1L2F_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2G_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2G_start : std_logic := '0';
  signal PC_L1L2G_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2HI_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2HI_start : std_logic := '0';
  signal PC_L1L2HI_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1L2JKL_bx : std_logic_vector(2 downto 0);
  signal PC_L1L2JKL_start : std_logic := '0';
  signal PC_L1L2JKL_bx_in : std_logic_vector(2 downto 0);
  signal PC_L2L3ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_L2L3ABCD_start : std_logic := '0';
  signal PC_L2L3ABCD_bx_in : std_logic_vector(2 downto 0);
  signal PC_L3L4AB_bx : std_logic_vector(2 downto 0);
  signal PC_L3L4AB_start : std_logic := '0';
  signal PC_L3L4AB_bx_in : std_logic_vector(2 downto 0);
  signal PC_L3L4CD_bx : std_logic_vector(2 downto 0);
  signal PC_L3L4CD_start : std_logic := '0';
  signal PC_L3L4CD_bx_in : std_logic_vector(2 downto 0);
  signal PC_L5L6ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_L5L6ABCD_start : std_logic := '0';
  signal PC_L5L6ABCD_bx_in : std_logic_vector(2 downto 0);
  signal PC_D1D2ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_D1D2ABCD_start : std_logic := '0';
  signal PC_D1D2ABCD_bx_in : std_logic_vector(2 downto 0);
  signal PC_D3D4ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_D3D4ABCD_start : std_logic := '0';
  signal PC_D3D4ABCD_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1D1ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_L1D1ABCD_start : std_logic := '0';
  signal PC_L1D1ABCD_bx_in : std_logic_vector(2 downto 0);
  signal PC_L1D1EFGH_bx : std_logic_vector(2 downto 0);
  signal PC_L1D1EFGH_start : std_logic := '0';
  signal PC_L1D1EFGH_bx_in : std_logic_vector(2 downto 0);
  signal PC_L2D1ABCD_bx : std_logic_vector(2 downto 0);
  signal PC_L2D1ABCD_start : std_logic := '0';
  signal PC_L2D1ABCD_bx_in : std_logic_vector(2 downto 0);
  signal VMSMER_done : std_logic := '0';
  signal VMSMER_bx_out : std_logic_vector(2 downto 0);
  signal VMSMER_bx_out_vld : std_logic;
  signal MP_L1PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIA_start : std_logic := '0';
  signal MP_L1PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIB_start : std_logic := '0';
  signal MP_L1PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIC_start : std_logic := '0';
  signal MP_L1PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHID_start : std_logic := '0';
  signal MP_L1PHIE_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIE_start : std_logic := '0';
  signal MP_L1PHIF_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIF_start : std_logic := '0';
  signal MP_L1PHIG_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIG_start : std_logic := '0';
  signal MP_L1PHIH_bx : std_logic_vector(2 downto 0);
  signal MP_L1PHIH_start : std_logic := '0';
  signal MP_L2PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L2PHIA_start : std_logic := '0';
  signal MP_L2PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L2PHIB_start : std_logic := '0';
  signal MP_L2PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L2PHIC_start : std_logic := '0';
  signal MP_L2PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L2PHID_start : std_logic := '0';
  signal MP_L3PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L3PHIA_start : std_logic := '0';
  signal MP_L3PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L3PHIB_start : std_logic := '0';
  signal MP_L3PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L3PHIC_start : std_logic := '0';
  signal MP_L3PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L3PHID_start : std_logic := '0';
  signal MP_L4PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L4PHIA_start : std_logic := '0';
  signal MP_L4PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L4PHIB_start : std_logic := '0';
  signal MP_L4PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L4PHIC_start : std_logic := '0';
  signal MP_L4PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L4PHID_start : std_logic := '0';
  signal MP_L5PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L5PHIA_start : std_logic := '0';
  signal MP_L5PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L5PHIB_start : std_logic := '0';
  signal MP_L5PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L5PHIC_start : std_logic := '0';
  signal MP_L5PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L5PHID_start : std_logic := '0';
  signal MP_L6PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_L6PHIA_start : std_logic := '0';
  signal MP_L6PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_L6PHIB_start : std_logic := '0';
  signal MP_L6PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_L6PHIC_start : std_logic := '0';
  signal MP_L6PHID_bx : std_logic_vector(2 downto 0);
  signal MP_L6PHID_start : std_logic := '0';
  signal MP_D1PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_D1PHIA_start : std_logic := '0';
  signal MP_D1PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_D1PHIB_start : std_logic := '0';
  signal MP_D1PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_D1PHIC_start : std_logic := '0';
  signal MP_D1PHID_bx : std_logic_vector(2 downto 0);
  signal MP_D1PHID_start : std_logic := '0';
  signal MP_D2PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_D2PHIA_start : std_logic := '0';
  signal MP_D2PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_D2PHIB_start : std_logic := '0';
  signal MP_D2PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_D2PHIC_start : std_logic := '0';
  signal MP_D2PHID_bx : std_logic_vector(2 downto 0);
  signal MP_D2PHID_start : std_logic := '0';
  signal MP_D3PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_D3PHIA_start : std_logic := '0';
  signal MP_D3PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_D3PHIB_start : std_logic := '0';
  signal MP_D3PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_D3PHIC_start : std_logic := '0';
  signal MP_D3PHID_bx : std_logic_vector(2 downto 0);
  signal MP_D3PHID_start : std_logic := '0';
  signal MP_D4PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_D4PHIA_start : std_logic := '0';
  signal MP_D4PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_D4PHIB_start : std_logic := '0';
  signal MP_D4PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_D4PHIC_start : std_logic := '0';
  signal MP_D4PHID_bx : std_logic_vector(2 downto 0);
  signal MP_D4PHID_start : std_logic := '0';
  signal MP_D5PHIA_bx : std_logic_vector(2 downto 0);
  signal MP_D5PHIA_start : std_logic := '0';
  signal MP_D5PHIB_bx : std_logic_vector(2 downto 0);
  signal MP_D5PHIB_start : std_logic := '0';
  signal MP_D5PHIC_bx : std_logic_vector(2 downto 0);
  signal MP_D5PHIC_start : std_logic := '0';
  signal MP_D5PHID_bx : std_logic_vector(2 downto 0);
  signal MP_D5PHID_start : std_logic := '0';
  signal MP_done : std_logic := '0';
  signal MP_bx_out : std_logic_vector(2 downto 0);
  signal MP_bx_out_vld : std_logic;
  signal TB_AAAA_bx : std_logic_vector(2 downto 0);
  signal TB_AAAA_start : std_logic := '0';
  signal TB_BBBB_bx : std_logic_vector(2 downto 0);
  signal TB_BBBB_start : std_logic := '0';

begin

    AS_L1PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIAin_wea_delay,
        addra     => AS_L1PHIAin_writeaddr_delay,
        dina      => AS_L1PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIAin_V_readaddr,
        doutb     => AS_L1PHIAin_V_dout,
        sync_nent => AS_L1PHIAin_start,
        nent_o    => AS_L1PHIAin_AV_dout_nent
      );

    AS_L1PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIAin_wea,
        addra     => AS_L1PHIAin_writeaddr,
        dina      => AS_L1PHIAin_din,
        wea_out       => AS_L1PHIAin_wea_delay,
        addra_out     => AS_L1PHIAin_writeaddr_delay,
        dina_out      => AS_L1PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIAin_start
      );

    AS_L1PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIBin_wea_delay,
        addra     => AS_L1PHIBin_writeaddr_delay,
        dina      => AS_L1PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIBin_V_readaddr,
        doutb     => AS_L1PHIBin_V_dout,
        sync_nent => AS_L1PHIBin_start,
        nent_o    => AS_L1PHIBin_AV_dout_nent
      );

    AS_L1PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIBin_wea,
        addra     => AS_L1PHIBin_writeaddr,
        dina      => AS_L1PHIBin_din,
        wea_out       => AS_L1PHIBin_wea_delay,
        addra_out     => AS_L1PHIBin_writeaddr_delay,
        dina_out      => AS_L1PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIBin_start
      );

    AS_L1PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHICin_wea_delay,
        addra     => AS_L1PHICin_writeaddr_delay,
        dina      => AS_L1PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHICin_V_readaddr,
        doutb     => AS_L1PHICin_V_dout,
        sync_nent => AS_L1PHICin_start,
        nent_o    => AS_L1PHICin_AV_dout_nent
      );

    AS_L1PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHICin_wea,
        addra     => AS_L1PHICin_writeaddr,
        dina      => AS_L1PHICin_din,
        wea_out       => AS_L1PHICin_wea_delay,
        addra_out     => AS_L1PHICin_writeaddr_delay,
        dina_out      => AS_L1PHICin_din_delay,
        done       => PC_start,
        start      => AS_L1PHICin_start
      );

    AS_L1PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIDin_wea_delay,
        addra     => AS_L1PHIDin_writeaddr_delay,
        dina      => AS_L1PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIDin_V_readaddr,
        doutb     => AS_L1PHIDin_V_dout,
        sync_nent => AS_L1PHIDin_start,
        nent_o    => AS_L1PHIDin_AV_dout_nent
      );

    AS_L1PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIDin_wea,
        addra     => AS_L1PHIDin_writeaddr,
        dina      => AS_L1PHIDin_din,
        wea_out       => AS_L1PHIDin_wea_delay,
        addra_out     => AS_L1PHIDin_writeaddr_delay,
        dina_out      => AS_L1PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIDin_start
      );

    AS_L1PHIEin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIEin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIEin_wea_delay,
        addra     => AS_L1PHIEin_writeaddr_delay,
        dina      => AS_L1PHIEin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIEin_V_readaddr,
        doutb     => AS_L1PHIEin_V_dout,
        sync_nent => AS_L1PHIEin_start,
        nent_o    => AS_L1PHIEin_AV_dout_nent
      );

    AS_L1PHIEin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIEin_wea,
        addra     => AS_L1PHIEin_writeaddr,
        dina      => AS_L1PHIEin_din,
        wea_out       => AS_L1PHIEin_wea_delay,
        addra_out     => AS_L1PHIEin_writeaddr_delay,
        dina_out      => AS_L1PHIEin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIEin_start
      );

    AS_L1PHIFin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIFin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIFin_wea_delay,
        addra     => AS_L1PHIFin_writeaddr_delay,
        dina      => AS_L1PHIFin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIFin_V_readaddr,
        doutb     => AS_L1PHIFin_V_dout,
        sync_nent => AS_L1PHIFin_start,
        nent_o    => AS_L1PHIFin_AV_dout_nent
      );

    AS_L1PHIFin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIFin_wea,
        addra     => AS_L1PHIFin_writeaddr,
        dina      => AS_L1PHIFin_din,
        wea_out       => AS_L1PHIFin_wea_delay,
        addra_out     => AS_L1PHIFin_writeaddr_delay,
        dina_out      => AS_L1PHIFin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIFin_start
      );

    AS_L1PHIGin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIGin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIGin_wea_delay,
        addra     => AS_L1PHIGin_writeaddr_delay,
        dina      => AS_L1PHIGin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIGin_V_readaddr,
        doutb     => AS_L1PHIGin_V_dout,
        sync_nent => AS_L1PHIGin_start,
        nent_o    => AS_L1PHIGin_AV_dout_nent
      );

    AS_L1PHIGin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIGin_wea,
        addra     => AS_L1PHIGin_writeaddr,
        dina      => AS_L1PHIGin_din,
        wea_out       => AS_L1PHIGin_wea_delay,
        addra_out     => AS_L1PHIGin_writeaddr_delay,
        dina_out      => AS_L1PHIGin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIGin_start
      );

    AS_L1PHIHin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIHin"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIHin_wea_delay,
        addra     => AS_L1PHIHin_writeaddr_delay,
        dina      => AS_L1PHIHin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIHin_V_readaddr,
        doutb     => AS_L1PHIHin_V_dout,
        sync_nent => AS_L1PHIHin_start,
        nent_o    => AS_L1PHIHin_AV_dout_nent
      );

    AS_L1PHIHin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIHin_wea,
        addra     => AS_L1PHIHin_writeaddr,
        dina      => AS_L1PHIHin_din,
        wea_out       => AS_L1PHIHin_wea_delay,
        addra_out     => AS_L1PHIHin_writeaddr_delay,
        dina_out      => AS_L1PHIHin_din_delay,
        done       => PC_start,
        start      => AS_L1PHIHin_start
      );

    AS_L2PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIAin_wea_delay,
        addra     => AS_L2PHIAin_writeaddr_delay,
        dina      => AS_L2PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIAin_V_readaddr,
        doutb     => AS_L2PHIAin_V_dout,
        sync_nent => AS_L2PHIAin_start,
        nent_o    => AS_L2PHIAin_AV_dout_nent
      );

    AS_L2PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIAin_wea,
        addra     => AS_L2PHIAin_writeaddr,
        dina      => AS_L2PHIAin_din,
        wea_out       => AS_L2PHIAin_wea_delay,
        addra_out     => AS_L2PHIAin_writeaddr_delay,
        dina_out      => AS_L2PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L2PHIAin_start
      );

    AS_L2PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIBin_wea_delay,
        addra     => AS_L2PHIBin_writeaddr_delay,
        dina      => AS_L2PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIBin_V_readaddr,
        doutb     => AS_L2PHIBin_V_dout,
        sync_nent => AS_L2PHIBin_start,
        nent_o    => AS_L2PHIBin_AV_dout_nent
      );

    AS_L2PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIBin_wea,
        addra     => AS_L2PHIBin_writeaddr,
        dina      => AS_L2PHIBin_din,
        wea_out       => AS_L2PHIBin_wea_delay,
        addra_out     => AS_L2PHIBin_writeaddr_delay,
        dina_out      => AS_L2PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L2PHIBin_start
      );

    AS_L2PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHICin_wea_delay,
        addra     => AS_L2PHICin_writeaddr_delay,
        dina      => AS_L2PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHICin_V_readaddr,
        doutb     => AS_L2PHICin_V_dout,
        sync_nent => AS_L2PHICin_start,
        nent_o    => AS_L2PHICin_AV_dout_nent
      );

    AS_L2PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHICin_wea,
        addra     => AS_L2PHICin_writeaddr,
        dina      => AS_L2PHICin_din,
        wea_out       => AS_L2PHICin_wea_delay,
        addra_out     => AS_L2PHICin_writeaddr_delay,
        dina_out      => AS_L2PHICin_din_delay,
        done       => PC_start,
        start      => AS_L2PHICin_start
      );

    AS_L2PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIDin_wea_delay,
        addra     => AS_L2PHIDin_writeaddr_delay,
        dina      => AS_L2PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIDin_V_readaddr,
        doutb     => AS_L2PHIDin_V_dout,
        sync_nent => AS_L2PHIDin_start,
        nent_o    => AS_L2PHIDin_AV_dout_nent
      );

    AS_L2PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIDin_wea,
        addra     => AS_L2PHIDin_writeaddr,
        dina      => AS_L2PHIDin_din,
        wea_out       => AS_L2PHIDin_wea_delay,
        addra_out     => AS_L2PHIDin_writeaddr_delay,
        dina_out      => AS_L2PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L2PHIDin_start
      );

    AS_L3PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIAin_wea_delay,
        addra     => AS_L3PHIAin_writeaddr_delay,
        dina      => AS_L3PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIAin_V_readaddr,
        doutb     => AS_L3PHIAin_V_dout,
        sync_nent => AS_L3PHIAin_start,
        nent_o    => AS_L3PHIAin_AV_dout_nent
      );

    AS_L3PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIAin_wea,
        addra     => AS_L3PHIAin_writeaddr,
        dina      => AS_L3PHIAin_din,
        wea_out       => AS_L3PHIAin_wea_delay,
        addra_out     => AS_L3PHIAin_writeaddr_delay,
        dina_out      => AS_L3PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L3PHIAin_start
      );

    AS_L3PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIBin_wea_delay,
        addra     => AS_L3PHIBin_writeaddr_delay,
        dina      => AS_L3PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIBin_V_readaddr,
        doutb     => AS_L3PHIBin_V_dout,
        sync_nent => AS_L3PHIBin_start,
        nent_o    => AS_L3PHIBin_AV_dout_nent
      );

    AS_L3PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIBin_wea,
        addra     => AS_L3PHIBin_writeaddr,
        dina      => AS_L3PHIBin_din,
        wea_out       => AS_L3PHIBin_wea_delay,
        addra_out     => AS_L3PHIBin_writeaddr_delay,
        dina_out      => AS_L3PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L3PHIBin_start
      );

    AS_L3PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHICin_wea_delay,
        addra     => AS_L3PHICin_writeaddr_delay,
        dina      => AS_L3PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHICin_V_readaddr,
        doutb     => AS_L3PHICin_V_dout,
        sync_nent => AS_L3PHICin_start,
        nent_o    => AS_L3PHICin_AV_dout_nent
      );

    AS_L3PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHICin_wea,
        addra     => AS_L3PHICin_writeaddr,
        dina      => AS_L3PHICin_din,
        wea_out       => AS_L3PHICin_wea_delay,
        addra_out     => AS_L3PHICin_writeaddr_delay,
        dina_out      => AS_L3PHICin_din_delay,
        done       => PC_start,
        start      => AS_L3PHICin_start
      );

    AS_L3PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIDin_wea_delay,
        addra     => AS_L3PHIDin_writeaddr_delay,
        dina      => AS_L3PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIDin_V_readaddr,
        doutb     => AS_L3PHIDin_V_dout,
        sync_nent => AS_L3PHIDin_start,
        nent_o    => AS_L3PHIDin_AV_dout_nent
      );

    AS_L3PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIDin_wea,
        addra     => AS_L3PHIDin_writeaddr,
        dina      => AS_L3PHIDin_din,
        wea_out       => AS_L3PHIDin_wea_delay,
        addra_out     => AS_L3PHIDin_writeaddr_delay,
        dina_out      => AS_L3PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L3PHIDin_start
      );

    AS_L4PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIAin_wea_delay,
        addra     => AS_L4PHIAin_writeaddr_delay,
        dina      => AS_L4PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIAin_V_readaddr,
        doutb     => AS_L4PHIAin_V_dout,
        sync_nent => AS_L4PHIAin_start,
        nent_o    => AS_L4PHIAin_AV_dout_nent
      );

    AS_L4PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIAin_wea,
        addra     => AS_L4PHIAin_writeaddr,
        dina      => AS_L4PHIAin_din,
        wea_out       => AS_L4PHIAin_wea_delay,
        addra_out     => AS_L4PHIAin_writeaddr_delay,
        dina_out      => AS_L4PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L4PHIAin_start
      );

    AS_L4PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIBin_wea_delay,
        addra     => AS_L4PHIBin_writeaddr_delay,
        dina      => AS_L4PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIBin_V_readaddr,
        doutb     => AS_L4PHIBin_V_dout,
        sync_nent => AS_L4PHIBin_start,
        nent_o    => AS_L4PHIBin_AV_dout_nent
      );

    AS_L4PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIBin_wea,
        addra     => AS_L4PHIBin_writeaddr,
        dina      => AS_L4PHIBin_din,
        wea_out       => AS_L4PHIBin_wea_delay,
        addra_out     => AS_L4PHIBin_writeaddr_delay,
        dina_out      => AS_L4PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L4PHIBin_start
      );

    AS_L4PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHICin_wea_delay,
        addra     => AS_L4PHICin_writeaddr_delay,
        dina      => AS_L4PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHICin_V_readaddr,
        doutb     => AS_L4PHICin_V_dout,
        sync_nent => AS_L4PHICin_start,
        nent_o    => AS_L4PHICin_AV_dout_nent
      );

    AS_L4PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHICin_wea,
        addra     => AS_L4PHICin_writeaddr,
        dina      => AS_L4PHICin_din,
        wea_out       => AS_L4PHICin_wea_delay,
        addra_out     => AS_L4PHICin_writeaddr_delay,
        dina_out      => AS_L4PHICin_din_delay,
        done       => PC_start,
        start      => AS_L4PHICin_start
      );

    AS_L4PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIDin_wea_delay,
        addra     => AS_L4PHIDin_writeaddr_delay,
        dina      => AS_L4PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIDin_V_readaddr,
        doutb     => AS_L4PHIDin_V_dout,
        sync_nent => AS_L4PHIDin_start,
        nent_o    => AS_L4PHIDin_AV_dout_nent
      );

    AS_L4PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIDin_wea,
        addra     => AS_L4PHIDin_writeaddr,
        dina      => AS_L4PHIDin_din,
        wea_out       => AS_L4PHIDin_wea_delay,
        addra_out     => AS_L4PHIDin_writeaddr_delay,
        dina_out      => AS_L4PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L4PHIDin_start
      );

    AS_L5PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIAin_wea_delay,
        addra     => AS_L5PHIAin_writeaddr_delay,
        dina      => AS_L5PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIAin_V_readaddr,
        doutb     => AS_L5PHIAin_V_dout,
        sync_nent => AS_L5PHIAin_start,
        nent_o    => AS_L5PHIAin_AV_dout_nent
      );

    AS_L5PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIAin_wea,
        addra     => AS_L5PHIAin_writeaddr,
        dina      => AS_L5PHIAin_din,
        wea_out       => AS_L5PHIAin_wea_delay,
        addra_out     => AS_L5PHIAin_writeaddr_delay,
        dina_out      => AS_L5PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L5PHIAin_start
      );

    AS_L5PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIBin_wea_delay,
        addra     => AS_L5PHIBin_writeaddr_delay,
        dina      => AS_L5PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIBin_V_readaddr,
        doutb     => AS_L5PHIBin_V_dout,
        sync_nent => AS_L5PHIBin_start,
        nent_o    => AS_L5PHIBin_AV_dout_nent
      );

    AS_L5PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIBin_wea,
        addra     => AS_L5PHIBin_writeaddr,
        dina      => AS_L5PHIBin_din,
        wea_out       => AS_L5PHIBin_wea_delay,
        addra_out     => AS_L5PHIBin_writeaddr_delay,
        dina_out      => AS_L5PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L5PHIBin_start
      );

    AS_L5PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHICin_wea_delay,
        addra     => AS_L5PHICin_writeaddr_delay,
        dina      => AS_L5PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHICin_V_readaddr,
        doutb     => AS_L5PHICin_V_dout,
        sync_nent => AS_L5PHICin_start,
        nent_o    => AS_L5PHICin_AV_dout_nent
      );

    AS_L5PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHICin_wea,
        addra     => AS_L5PHICin_writeaddr,
        dina      => AS_L5PHICin_din,
        wea_out       => AS_L5PHICin_wea_delay,
        addra_out     => AS_L5PHICin_writeaddr_delay,
        dina_out      => AS_L5PHICin_din_delay,
        done       => PC_start,
        start      => AS_L5PHICin_start
      );

    AS_L5PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIDin_wea_delay,
        addra     => AS_L5PHIDin_writeaddr_delay,
        dina      => AS_L5PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIDin_V_readaddr,
        doutb     => AS_L5PHIDin_V_dout,
        sync_nent => AS_L5PHIDin_start,
        nent_o    => AS_L5PHIDin_AV_dout_nent
      );

    AS_L5PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIDin_wea,
        addra     => AS_L5PHIDin_writeaddr,
        dina      => AS_L5PHIDin_din,
        wea_out       => AS_L5PHIDin_wea_delay,
        addra_out     => AS_L5PHIDin_writeaddr_delay,
        dina_out      => AS_L5PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L5PHIDin_start
      );

    AS_L6PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIAin_wea_delay,
        addra     => AS_L6PHIAin_writeaddr_delay,
        dina      => AS_L6PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIAin_V_readaddr,
        doutb     => AS_L6PHIAin_V_dout,
        sync_nent => AS_L6PHIAin_start,
        nent_o    => AS_L6PHIAin_AV_dout_nent
      );

    AS_L6PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIAin_wea,
        addra     => AS_L6PHIAin_writeaddr,
        dina      => AS_L6PHIAin_din,
        wea_out       => AS_L6PHIAin_wea_delay,
        addra_out     => AS_L6PHIAin_writeaddr_delay,
        dina_out      => AS_L6PHIAin_din_delay,
        done       => PC_start,
        start      => AS_L6PHIAin_start
      );

    AS_L6PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIBin_wea_delay,
        addra     => AS_L6PHIBin_writeaddr_delay,
        dina      => AS_L6PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIBin_V_readaddr,
        doutb     => AS_L6PHIBin_V_dout,
        sync_nent => AS_L6PHIBin_start,
        nent_o    => AS_L6PHIBin_AV_dout_nent
      );

    AS_L6PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIBin_wea,
        addra     => AS_L6PHIBin_writeaddr,
        dina      => AS_L6PHIBin_din,
        wea_out       => AS_L6PHIBin_wea_delay,
        addra_out     => AS_L6PHIBin_writeaddr_delay,
        dina_out      => AS_L6PHIBin_din_delay,
        done       => PC_start,
        start      => AS_L6PHIBin_start
      );

    AS_L6PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHICin_wea_delay,
        addra     => AS_L6PHICin_writeaddr_delay,
        dina      => AS_L6PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHICin_V_readaddr,
        doutb     => AS_L6PHICin_V_dout,
        sync_nent => AS_L6PHICin_start,
        nent_o    => AS_L6PHICin_AV_dout_nent
      );

    AS_L6PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHICin_wea,
        addra     => AS_L6PHICin_writeaddr,
        dina      => AS_L6PHICin_din,
        wea_out       => AS_L6PHICin_wea_delay,
        addra_out     => AS_L6PHICin_writeaddr_delay,
        dina_out      => AS_L6PHICin_din_delay,
        done       => PC_start,
        start      => AS_L6PHICin_start
      );

    AS_L6PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIDin_wea_delay,
        addra     => AS_L6PHIDin_writeaddr_delay,
        dina      => AS_L6PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIDin_V_readaddr,
        doutb     => AS_L6PHIDin_V_dout,
        sync_nent => AS_L6PHIDin_start,
        nent_o    => AS_L6PHIDin_AV_dout_nent
      );

    AS_L6PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIDin_wea,
        addra     => AS_L6PHIDin_writeaddr,
        dina      => AS_L6PHIDin_din,
        wea_out       => AS_L6PHIDin_wea_delay,
        addra_out     => AS_L6PHIDin_writeaddr_delay,
        dina_out      => AS_L6PHIDin_din_delay,
        done       => PC_start,
        start      => AS_L6PHIDin_start
      );

    AS_D1PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIAin_wea_delay,
        addra     => AS_D1PHIAin_writeaddr_delay,
        dina      => AS_D1PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIAin_V_readaddr,
        doutb     => AS_D1PHIAin_V_dout,
        sync_nent => AS_D1PHIAin_start,
        nent_o    => AS_D1PHIAin_AV_dout_nent
      );

    AS_D1PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIAin_wea,
        addra     => AS_D1PHIAin_writeaddr,
        dina      => AS_D1PHIAin_din,
        wea_out       => AS_D1PHIAin_wea_delay,
        addra_out     => AS_D1PHIAin_writeaddr_delay,
        dina_out      => AS_D1PHIAin_din_delay,
        done       => PC_start,
        start      => AS_D1PHIAin_start
      );

    AS_D1PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIBin_wea_delay,
        addra     => AS_D1PHIBin_writeaddr_delay,
        dina      => AS_D1PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIBin_V_readaddr,
        doutb     => AS_D1PHIBin_V_dout,
        sync_nent => AS_D1PHIBin_start,
        nent_o    => AS_D1PHIBin_AV_dout_nent
      );

    AS_D1PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIBin_wea,
        addra     => AS_D1PHIBin_writeaddr,
        dina      => AS_D1PHIBin_din,
        wea_out       => AS_D1PHIBin_wea_delay,
        addra_out     => AS_D1PHIBin_writeaddr_delay,
        dina_out      => AS_D1PHIBin_din_delay,
        done       => PC_start,
        start      => AS_D1PHIBin_start
      );

    AS_D1PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHICin_wea_delay,
        addra     => AS_D1PHICin_writeaddr_delay,
        dina      => AS_D1PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHICin_V_readaddr,
        doutb     => AS_D1PHICin_V_dout,
        sync_nent => AS_D1PHICin_start,
        nent_o    => AS_D1PHICin_AV_dout_nent
      );

    AS_D1PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHICin_wea,
        addra     => AS_D1PHICin_writeaddr,
        dina      => AS_D1PHICin_din,
        wea_out       => AS_D1PHICin_wea_delay,
        addra_out     => AS_D1PHICin_writeaddr_delay,
        dina_out      => AS_D1PHICin_din_delay,
        done       => PC_start,
        start      => AS_D1PHICin_start
      );

    AS_D1PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIDin_wea_delay,
        addra     => AS_D1PHIDin_writeaddr_delay,
        dina      => AS_D1PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIDin_V_readaddr,
        doutb     => AS_D1PHIDin_V_dout,
        sync_nent => AS_D1PHIDin_start,
        nent_o    => AS_D1PHIDin_AV_dout_nent
      );

    AS_D1PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIDin_wea,
        addra     => AS_D1PHIDin_writeaddr,
        dina      => AS_D1PHIDin_din,
        wea_out       => AS_D1PHIDin_wea_delay,
        addra_out     => AS_D1PHIDin_writeaddr_delay,
        dina_out      => AS_D1PHIDin_din_delay,
        done       => PC_start,
        start      => AS_D1PHIDin_start
      );

    AS_D2PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIAin_wea_delay,
        addra     => AS_D2PHIAin_writeaddr_delay,
        dina      => AS_D2PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIAin_V_readaddr,
        doutb     => AS_D2PHIAin_V_dout,
        sync_nent => AS_D2PHIAin_start,
        nent_o    => AS_D2PHIAin_AV_dout_nent
      );

    AS_D2PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIAin_wea,
        addra     => AS_D2PHIAin_writeaddr,
        dina      => AS_D2PHIAin_din,
        wea_out       => AS_D2PHIAin_wea_delay,
        addra_out     => AS_D2PHIAin_writeaddr_delay,
        dina_out      => AS_D2PHIAin_din_delay,
        done       => PC_start,
        start      => AS_D2PHIAin_start
      );

    AS_D2PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIBin_wea_delay,
        addra     => AS_D2PHIBin_writeaddr_delay,
        dina      => AS_D2PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIBin_V_readaddr,
        doutb     => AS_D2PHIBin_V_dout,
        sync_nent => AS_D2PHIBin_start,
        nent_o    => AS_D2PHIBin_AV_dout_nent
      );

    AS_D2PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIBin_wea,
        addra     => AS_D2PHIBin_writeaddr,
        dina      => AS_D2PHIBin_din,
        wea_out       => AS_D2PHIBin_wea_delay,
        addra_out     => AS_D2PHIBin_writeaddr_delay,
        dina_out      => AS_D2PHIBin_din_delay,
        done       => PC_start,
        start      => AS_D2PHIBin_start
      );

    AS_D2PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHICin_wea_delay,
        addra     => AS_D2PHICin_writeaddr_delay,
        dina      => AS_D2PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHICin_V_readaddr,
        doutb     => AS_D2PHICin_V_dout,
        sync_nent => AS_D2PHICin_start,
        nent_o    => AS_D2PHICin_AV_dout_nent
      );

    AS_D2PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHICin_wea,
        addra     => AS_D2PHICin_writeaddr,
        dina      => AS_D2PHICin_din,
        wea_out       => AS_D2PHICin_wea_delay,
        addra_out     => AS_D2PHICin_writeaddr_delay,
        dina_out      => AS_D2PHICin_din_delay,
        done       => PC_start,
        start      => AS_D2PHICin_start
      );

    AS_D2PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIDin_wea_delay,
        addra     => AS_D2PHIDin_writeaddr_delay,
        dina      => AS_D2PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIDin_V_readaddr,
        doutb     => AS_D2PHIDin_V_dout,
        sync_nent => AS_D2PHIDin_start,
        nent_o    => AS_D2PHIDin_AV_dout_nent
      );

    AS_D2PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIDin_wea,
        addra     => AS_D2PHIDin_writeaddr,
        dina      => AS_D2PHIDin_din,
        wea_out       => AS_D2PHIDin_wea_delay,
        addra_out     => AS_D2PHIDin_writeaddr_delay,
        dina_out      => AS_D2PHIDin_din_delay,
        done       => PC_start,
        start      => AS_D2PHIDin_start
      );

    AS_D3PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIAin_wea_delay,
        addra     => AS_D3PHIAin_writeaddr_delay,
        dina      => AS_D3PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIAin_V_readaddr,
        doutb     => AS_D3PHIAin_V_dout,
        sync_nent => AS_D3PHIAin_start,
        nent_o    => AS_D3PHIAin_AV_dout_nent
      );

    AS_D3PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIAin_wea,
        addra     => AS_D3PHIAin_writeaddr,
        dina      => AS_D3PHIAin_din,
        wea_out       => AS_D3PHIAin_wea_delay,
        addra_out     => AS_D3PHIAin_writeaddr_delay,
        dina_out      => AS_D3PHIAin_din_delay,
        done       => PC_start,
        start      => AS_D3PHIAin_start
      );

    AS_D3PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIBin_wea_delay,
        addra     => AS_D3PHIBin_writeaddr_delay,
        dina      => AS_D3PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIBin_V_readaddr,
        doutb     => AS_D3PHIBin_V_dout,
        sync_nent => AS_D3PHIBin_start,
        nent_o    => AS_D3PHIBin_AV_dout_nent
      );

    AS_D3PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIBin_wea,
        addra     => AS_D3PHIBin_writeaddr,
        dina      => AS_D3PHIBin_din,
        wea_out       => AS_D3PHIBin_wea_delay,
        addra_out     => AS_D3PHIBin_writeaddr_delay,
        dina_out      => AS_D3PHIBin_din_delay,
        done       => PC_start,
        start      => AS_D3PHIBin_start
      );

    AS_D3PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHICin_wea_delay,
        addra     => AS_D3PHICin_writeaddr_delay,
        dina      => AS_D3PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHICin_V_readaddr,
        doutb     => AS_D3PHICin_V_dout,
        sync_nent => AS_D3PHICin_start,
        nent_o    => AS_D3PHICin_AV_dout_nent
      );

    AS_D3PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHICin_wea,
        addra     => AS_D3PHICin_writeaddr,
        dina      => AS_D3PHICin_din,
        wea_out       => AS_D3PHICin_wea_delay,
        addra_out     => AS_D3PHICin_writeaddr_delay,
        dina_out      => AS_D3PHICin_din_delay,
        done       => PC_start,
        start      => AS_D3PHICin_start
      );

    AS_D3PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIDin_wea_delay,
        addra     => AS_D3PHIDin_writeaddr_delay,
        dina      => AS_D3PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIDin_V_readaddr,
        doutb     => AS_D3PHIDin_V_dout,
        sync_nent => AS_D3PHIDin_start,
        nent_o    => AS_D3PHIDin_AV_dout_nent
      );

    AS_D3PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIDin_wea,
        addra     => AS_D3PHIDin_writeaddr,
        dina      => AS_D3PHIDin_din,
        wea_out       => AS_D3PHIDin_wea_delay,
        addra_out     => AS_D3PHIDin_writeaddr_delay,
        dina_out      => AS_D3PHIDin_din_delay,
        done       => PC_start,
        start      => AS_D3PHIDin_start
      );

    AS_D4PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIAin_wea_delay,
        addra     => AS_D4PHIAin_writeaddr_delay,
        dina      => AS_D4PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIAin_V_readaddr,
        doutb     => AS_D4PHIAin_V_dout,
        sync_nent => AS_D4PHIAin_start,
        nent_o    => AS_D4PHIAin_AV_dout_nent
      );

    AS_D4PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIAin_wea,
        addra     => AS_D4PHIAin_writeaddr,
        dina      => AS_D4PHIAin_din,
        wea_out       => AS_D4PHIAin_wea_delay,
        addra_out     => AS_D4PHIAin_writeaddr_delay,
        dina_out      => AS_D4PHIAin_din_delay,
        done       => PC_start,
        start      => AS_D4PHIAin_start
      );

    AS_D4PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIBin_wea_delay,
        addra     => AS_D4PHIBin_writeaddr_delay,
        dina      => AS_D4PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIBin_V_readaddr,
        doutb     => AS_D4PHIBin_V_dout,
        sync_nent => AS_D4PHIBin_start,
        nent_o    => AS_D4PHIBin_AV_dout_nent
      );

    AS_D4PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIBin_wea,
        addra     => AS_D4PHIBin_writeaddr,
        dina      => AS_D4PHIBin_din,
        wea_out       => AS_D4PHIBin_wea_delay,
        addra_out     => AS_D4PHIBin_writeaddr_delay,
        dina_out      => AS_D4PHIBin_din_delay,
        done       => PC_start,
        start      => AS_D4PHIBin_start
      );

    AS_D4PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHICin_wea_delay,
        addra     => AS_D4PHICin_writeaddr_delay,
        dina      => AS_D4PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHICin_V_readaddr,
        doutb     => AS_D4PHICin_V_dout,
        sync_nent => AS_D4PHICin_start,
        nent_o    => AS_D4PHICin_AV_dout_nent
      );

    AS_D4PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHICin_wea,
        addra     => AS_D4PHICin_writeaddr,
        dina      => AS_D4PHICin_din,
        wea_out       => AS_D4PHICin_wea_delay,
        addra_out     => AS_D4PHICin_writeaddr_delay,
        dina_out      => AS_D4PHICin_din_delay,
        done       => PC_start,
        start      => AS_D4PHICin_start
      );

    AS_D4PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIDin_wea_delay,
        addra     => AS_D4PHIDin_writeaddr_delay,
        dina      => AS_D4PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIDin_V_readaddr,
        doutb     => AS_D4PHIDin_V_dout,
        sync_nent => AS_D4PHIDin_start,
        nent_o    => AS_D4PHIDin_AV_dout_nent
      );

    AS_D4PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIDin_wea,
        addra     => AS_D4PHIDin_writeaddr,
        dina      => AS_D4PHIDin_din,
        wea_out       => AS_D4PHIDin_wea_delay,
        addra_out     => AS_D4PHIDin_writeaddr_delay,
        dina_out      => AS_D4PHIDin_din_delay,
        done       => PC_start,
        start      => AS_D4PHIDin_start
      );

    AS_D5PHIAin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIAin"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIAin_wea_delay,
        addra     => AS_D5PHIAin_writeaddr_delay,
        dina      => AS_D5PHIAin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIAin_V_readaddr,
        doutb     => AS_D5PHIAin_V_dout,
        sync_nent => AS_D5PHIAin_start,
        nent_o    => AS_D5PHIAin_AV_dout_nent
      );

    AS_D5PHIAin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIAin_wea,
        addra     => AS_D5PHIAin_writeaddr,
        dina      => AS_D5PHIAin_din,
        wea_out       => AS_D5PHIAin_wea_delay,
        addra_out     => AS_D5PHIAin_writeaddr_delay,
        dina_out      => AS_D5PHIAin_din_delay,
        done       => PC_start,
        start      => AS_D5PHIAin_start
      );

    AS_D5PHIBin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIBin"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIBin_wea_delay,
        addra     => AS_D5PHIBin_writeaddr_delay,
        dina      => AS_D5PHIBin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIBin_V_readaddr,
        doutb     => AS_D5PHIBin_V_dout,
        sync_nent => AS_D5PHIBin_start,
        nent_o    => AS_D5PHIBin_AV_dout_nent
      );

    AS_D5PHIBin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIBin_wea,
        addra     => AS_D5PHIBin_writeaddr,
        dina      => AS_D5PHIBin_din,
        wea_out       => AS_D5PHIBin_wea_delay,
        addra_out     => AS_D5PHIBin_writeaddr_delay,
        dina_out      => AS_D5PHIBin_din_delay,
        done       => PC_start,
        start      => AS_D5PHIBin_start
      );

    AS_D5PHICin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHICin"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHICin_wea_delay,
        addra     => AS_D5PHICin_writeaddr_delay,
        dina      => AS_D5PHICin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHICin_V_readaddr,
        doutb     => AS_D5PHICin_V_dout,
        sync_nent => AS_D5PHICin_start,
        nent_o    => AS_D5PHICin_AV_dout_nent
      );

    AS_D5PHICin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHICin_wea,
        addra     => AS_D5PHICin_writeaddr,
        dina      => AS_D5PHICin_din,
        wea_out       => AS_D5PHICin_wea_delay,
        addra_out     => AS_D5PHICin_writeaddr_delay,
        dina_out      => AS_D5PHICin_din_delay,
        done       => PC_start,
        start      => AS_D5PHICin_start
      );

    AS_D5PHIDin : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIDin"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIDin_wea_delay,
        addra     => AS_D5PHIDin_writeaddr_delay,
        dina      => AS_D5PHIDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIDin_V_readaddr,
        doutb     => AS_D5PHIDin_V_dout,
        sync_nent => AS_D5PHIDin_start,
        nent_o    => AS_D5PHIDin_AV_dout_nent
      );

    AS_D5PHIDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIDin_wea,
        addra     => AS_D5PHIDin_writeaddr,
        dina      => AS_D5PHIDin_din,
        wea_out       => AS_D5PHIDin_wea_delay,
        addra_out     => AS_D5PHIDin_writeaddr_delay,
        dina_out      => AS_D5PHIDin_din_delay,
        done       => PC_start,
        start      => AS_D5PHIDin_start
      );

    AS_L1PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIAn2_wea_delay,
        addra     => AS_L1PHIAn2_writeaddr_delay,
        dina      => AS_L1PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIAn2_V_readaddr,
        doutb     => AS_L1PHIAn2_V_dout,
        sync_nent => AS_L1PHIAn2_start,
        nent_o    => open
      );

    AS_L1PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIAn2_wea,
        addra     => AS_L1PHIAn2_writeaddr,
        dina      => AS_L1PHIAn2_din,
        wea_out       => AS_L1PHIAn2_wea_delay,
        addra_out     => AS_L1PHIAn2_writeaddr_delay,
        dina_out      => AS_L1PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIAn2_start
      );

    AS_L1PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIBn2_wea_delay,
        addra     => AS_L1PHIBn2_writeaddr_delay,
        dina      => AS_L1PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIBn2_V_readaddr,
        doutb     => AS_L1PHIBn2_V_dout,
        sync_nent => AS_L1PHIBn2_start,
        nent_o    => open
      );

    AS_L1PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIBn2_wea,
        addra     => AS_L1PHIBn2_writeaddr,
        dina      => AS_L1PHIBn2_din,
        wea_out       => AS_L1PHIBn2_wea_delay,
        addra_out     => AS_L1PHIBn2_writeaddr_delay,
        dina_out      => AS_L1PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIBn2_start
      );

    AS_L1PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHICn2_wea_delay,
        addra     => AS_L1PHICn2_writeaddr_delay,
        dina      => AS_L1PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHICn2_V_readaddr,
        doutb     => AS_L1PHICn2_V_dout,
        sync_nent => AS_L1PHICn2_start,
        nent_o    => open
      );

    AS_L1PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHICn2_wea,
        addra     => AS_L1PHICn2_writeaddr,
        dina      => AS_L1PHICn2_din,
        wea_out       => AS_L1PHICn2_wea_delay,
        addra_out     => AS_L1PHICn2_writeaddr_delay,
        dina_out      => AS_L1PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHICn2_start
      );

    AS_L1PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIDn2_wea_delay,
        addra     => AS_L1PHIDn2_writeaddr_delay,
        dina      => AS_L1PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIDn2_V_readaddr,
        doutb     => AS_L1PHIDn2_V_dout,
        sync_nent => AS_L1PHIDn2_start,
        nent_o    => open
      );

    AS_L1PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIDn2_wea,
        addra     => AS_L1PHIDn2_writeaddr,
        dina      => AS_L1PHIDn2_din,
        wea_out       => AS_L1PHIDn2_wea_delay,
        addra_out     => AS_L1PHIDn2_writeaddr_delay,
        dina_out      => AS_L1PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIDn2_start
      );

    AS_L1PHIEn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIEn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIEn2_wea_delay,
        addra     => AS_L1PHIEn2_writeaddr_delay,
        dina      => AS_L1PHIEn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIEn2_V_readaddr,
        doutb     => AS_L1PHIEn2_V_dout,
        sync_nent => AS_L1PHIEn2_start,
        nent_o    => open
      );

    AS_L1PHIEn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIEn2_wea,
        addra     => AS_L1PHIEn2_writeaddr,
        dina      => AS_L1PHIEn2_din,
        wea_out       => AS_L1PHIEn2_wea_delay,
        addra_out     => AS_L1PHIEn2_writeaddr_delay,
        dina_out      => AS_L1PHIEn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIEn2_start
      );

    AS_L1PHIFn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIFn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIFn2_wea_delay,
        addra     => AS_L1PHIFn2_writeaddr_delay,
        dina      => AS_L1PHIFn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIFn2_V_readaddr,
        doutb     => AS_L1PHIFn2_V_dout,
        sync_nent => AS_L1PHIFn2_start,
        nent_o    => open
      );

    AS_L1PHIFn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIFn2_wea,
        addra     => AS_L1PHIFn2_writeaddr,
        dina      => AS_L1PHIFn2_din,
        wea_out       => AS_L1PHIFn2_wea_delay,
        addra_out     => AS_L1PHIFn2_writeaddr_delay,
        dina_out      => AS_L1PHIFn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIFn2_start
      );

    AS_L1PHIGn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIGn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIGn2_wea_delay,
        addra     => AS_L1PHIGn2_writeaddr_delay,
        dina      => AS_L1PHIGn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIGn2_V_readaddr,
        doutb     => AS_L1PHIGn2_V_dout,
        sync_nent => AS_L1PHIGn2_start,
        nent_o    => open
      );

    AS_L1PHIGn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIGn2_wea,
        addra     => AS_L1PHIGn2_writeaddr,
        dina      => AS_L1PHIGn2_din,
        wea_out       => AS_L1PHIGn2_wea_delay,
        addra_out     => AS_L1PHIGn2_writeaddr_delay,
        dina_out      => AS_L1PHIGn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIGn2_start
      );

    AS_L1PHIHn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIHn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIHn2_wea_delay,
        addra     => AS_L1PHIHn2_writeaddr_delay,
        dina      => AS_L1PHIHn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIHn2_V_readaddr,
        doutb     => AS_L1PHIHn2_V_dout,
        sync_nent => AS_L1PHIHn2_start,
        nent_o    => open
      );

    AS_L1PHIHn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIHn2_wea,
        addra     => AS_L1PHIHn2_writeaddr,
        dina      => AS_L1PHIHn2_din,
        wea_out       => AS_L1PHIHn2_wea_delay,
        addra_out     => AS_L1PHIHn2_writeaddr_delay,
        dina_out      => AS_L1PHIHn2_din_delay,
        done       => PC_done,
        start      => AS_L1PHIHn2_start
      );

    AS_L2PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIAn2_wea_delay,
        addra     => AS_L2PHIAn2_writeaddr_delay,
        dina      => AS_L2PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIAn2_V_readaddr,
        doutb     => AS_L2PHIAn2_V_dout,
        sync_nent => AS_L2PHIAn2_start,
        nent_o    => open
      );

    AS_L2PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIAn2_wea,
        addra     => AS_L2PHIAn2_writeaddr,
        dina      => AS_L2PHIAn2_din,
        wea_out       => AS_L2PHIAn2_wea_delay,
        addra_out     => AS_L2PHIAn2_writeaddr_delay,
        dina_out      => AS_L2PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L2PHIAn2_start
      );

    AS_L2PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIBn2_wea_delay,
        addra     => AS_L2PHIBn2_writeaddr_delay,
        dina      => AS_L2PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIBn2_V_readaddr,
        doutb     => AS_L2PHIBn2_V_dout,
        sync_nent => AS_L2PHIBn2_start,
        nent_o    => open
      );

    AS_L2PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIBn2_wea,
        addra     => AS_L2PHIBn2_writeaddr,
        dina      => AS_L2PHIBn2_din,
        wea_out       => AS_L2PHIBn2_wea_delay,
        addra_out     => AS_L2PHIBn2_writeaddr_delay,
        dina_out      => AS_L2PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L2PHIBn2_start
      );

    AS_L2PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHICn2_wea_delay,
        addra     => AS_L2PHICn2_writeaddr_delay,
        dina      => AS_L2PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHICn2_V_readaddr,
        doutb     => AS_L2PHICn2_V_dout,
        sync_nent => AS_L2PHICn2_start,
        nent_o    => open
      );

    AS_L2PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHICn2_wea,
        addra     => AS_L2PHICn2_writeaddr,
        dina      => AS_L2PHICn2_din,
        wea_out       => AS_L2PHICn2_wea_delay,
        addra_out     => AS_L2PHICn2_writeaddr_delay,
        dina_out      => AS_L2PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L2PHICn2_start
      );

    AS_L2PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIDn2_wea_delay,
        addra     => AS_L2PHIDn2_writeaddr_delay,
        dina      => AS_L2PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIDn2_V_readaddr,
        doutb     => AS_L2PHIDn2_V_dout,
        sync_nent => AS_L2PHIDn2_start,
        nent_o    => open
      );

    AS_L2PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIDn2_wea,
        addra     => AS_L2PHIDn2_writeaddr,
        dina      => AS_L2PHIDn2_din,
        wea_out       => AS_L2PHIDn2_wea_delay,
        addra_out     => AS_L2PHIDn2_writeaddr_delay,
        dina_out      => AS_L2PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L2PHIDn2_start
      );

    AS_L3PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIAn2_wea_delay,
        addra     => AS_L3PHIAn2_writeaddr_delay,
        dina      => AS_L3PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIAn2_V_readaddr,
        doutb     => AS_L3PHIAn2_V_dout,
        sync_nent => AS_L3PHIAn2_start,
        nent_o    => open
      );

    AS_L3PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIAn2_wea,
        addra     => AS_L3PHIAn2_writeaddr,
        dina      => AS_L3PHIAn2_din,
        wea_out       => AS_L3PHIAn2_wea_delay,
        addra_out     => AS_L3PHIAn2_writeaddr_delay,
        dina_out      => AS_L3PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L3PHIAn2_start
      );

    AS_L3PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIBn2_wea_delay,
        addra     => AS_L3PHIBn2_writeaddr_delay,
        dina      => AS_L3PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIBn2_V_readaddr,
        doutb     => AS_L3PHIBn2_V_dout,
        sync_nent => AS_L3PHIBn2_start,
        nent_o    => open
      );

    AS_L3PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIBn2_wea,
        addra     => AS_L3PHIBn2_writeaddr,
        dina      => AS_L3PHIBn2_din,
        wea_out       => AS_L3PHIBn2_wea_delay,
        addra_out     => AS_L3PHIBn2_writeaddr_delay,
        dina_out      => AS_L3PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L3PHIBn2_start
      );

    AS_L3PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHICn2_wea_delay,
        addra     => AS_L3PHICn2_writeaddr_delay,
        dina      => AS_L3PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHICn2_V_readaddr,
        doutb     => AS_L3PHICn2_V_dout,
        sync_nent => AS_L3PHICn2_start,
        nent_o    => open
      );

    AS_L3PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHICn2_wea,
        addra     => AS_L3PHICn2_writeaddr,
        dina      => AS_L3PHICn2_din,
        wea_out       => AS_L3PHICn2_wea_delay,
        addra_out     => AS_L3PHICn2_writeaddr_delay,
        dina_out      => AS_L3PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L3PHICn2_start
      );

    AS_L3PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIDn2_wea_delay,
        addra     => AS_L3PHIDn2_writeaddr_delay,
        dina      => AS_L3PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIDn2_V_readaddr,
        doutb     => AS_L3PHIDn2_V_dout,
        sync_nent => AS_L3PHIDn2_start,
        nent_o    => open
      );

    AS_L3PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIDn2_wea,
        addra     => AS_L3PHIDn2_writeaddr,
        dina      => AS_L3PHIDn2_din,
        wea_out       => AS_L3PHIDn2_wea_delay,
        addra_out     => AS_L3PHIDn2_writeaddr_delay,
        dina_out      => AS_L3PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L3PHIDn2_start
      );

    AS_L4PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIAn2_wea_delay,
        addra     => AS_L4PHIAn2_writeaddr_delay,
        dina      => AS_L4PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIAn2_V_readaddr,
        doutb     => AS_L4PHIAn2_V_dout,
        sync_nent => AS_L4PHIAn2_start,
        nent_o    => open
      );

    AS_L4PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIAn2_wea,
        addra     => AS_L4PHIAn2_writeaddr,
        dina      => AS_L4PHIAn2_din,
        wea_out       => AS_L4PHIAn2_wea_delay,
        addra_out     => AS_L4PHIAn2_writeaddr_delay,
        dina_out      => AS_L4PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L4PHIAn2_start
      );

    AS_L4PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIBn2_wea_delay,
        addra     => AS_L4PHIBn2_writeaddr_delay,
        dina      => AS_L4PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIBn2_V_readaddr,
        doutb     => AS_L4PHIBn2_V_dout,
        sync_nent => AS_L4PHIBn2_start,
        nent_o    => open
      );

    AS_L4PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIBn2_wea,
        addra     => AS_L4PHIBn2_writeaddr,
        dina      => AS_L4PHIBn2_din,
        wea_out       => AS_L4PHIBn2_wea_delay,
        addra_out     => AS_L4PHIBn2_writeaddr_delay,
        dina_out      => AS_L4PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L4PHIBn2_start
      );

    AS_L4PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHICn2_wea_delay,
        addra     => AS_L4PHICn2_writeaddr_delay,
        dina      => AS_L4PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHICn2_V_readaddr,
        doutb     => AS_L4PHICn2_V_dout,
        sync_nent => AS_L4PHICn2_start,
        nent_o    => open
      );

    AS_L4PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHICn2_wea,
        addra     => AS_L4PHICn2_writeaddr,
        dina      => AS_L4PHICn2_din,
        wea_out       => AS_L4PHICn2_wea_delay,
        addra_out     => AS_L4PHICn2_writeaddr_delay,
        dina_out      => AS_L4PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L4PHICn2_start
      );

    AS_L4PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIDn2_wea_delay,
        addra     => AS_L4PHIDn2_writeaddr_delay,
        dina      => AS_L4PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIDn2_V_readaddr,
        doutb     => AS_L4PHIDn2_V_dout,
        sync_nent => AS_L4PHIDn2_start,
        nent_o    => open
      );

    AS_L4PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIDn2_wea,
        addra     => AS_L4PHIDn2_writeaddr,
        dina      => AS_L4PHIDn2_din,
        wea_out       => AS_L4PHIDn2_wea_delay,
        addra_out     => AS_L4PHIDn2_writeaddr_delay,
        dina_out      => AS_L4PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L4PHIDn2_start
      );

    AS_L5PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIAn2_wea_delay,
        addra     => AS_L5PHIAn2_writeaddr_delay,
        dina      => AS_L5PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIAn2_V_readaddr,
        doutb     => AS_L5PHIAn2_V_dout,
        sync_nent => AS_L5PHIAn2_start,
        nent_o    => open
      );

    AS_L5PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIAn2_wea,
        addra     => AS_L5PHIAn2_writeaddr,
        dina      => AS_L5PHIAn2_din,
        wea_out       => AS_L5PHIAn2_wea_delay,
        addra_out     => AS_L5PHIAn2_writeaddr_delay,
        dina_out      => AS_L5PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L5PHIAn2_start
      );

    AS_L5PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIBn2_wea_delay,
        addra     => AS_L5PHIBn2_writeaddr_delay,
        dina      => AS_L5PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIBn2_V_readaddr,
        doutb     => AS_L5PHIBn2_V_dout,
        sync_nent => AS_L5PHIBn2_start,
        nent_o    => open
      );

    AS_L5PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIBn2_wea,
        addra     => AS_L5PHIBn2_writeaddr,
        dina      => AS_L5PHIBn2_din,
        wea_out       => AS_L5PHIBn2_wea_delay,
        addra_out     => AS_L5PHIBn2_writeaddr_delay,
        dina_out      => AS_L5PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L5PHIBn2_start
      );

    AS_L5PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHICn2_wea_delay,
        addra     => AS_L5PHICn2_writeaddr_delay,
        dina      => AS_L5PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHICn2_V_readaddr,
        doutb     => AS_L5PHICn2_V_dout,
        sync_nent => AS_L5PHICn2_start,
        nent_o    => open
      );

    AS_L5PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHICn2_wea,
        addra     => AS_L5PHICn2_writeaddr,
        dina      => AS_L5PHICn2_din,
        wea_out       => AS_L5PHICn2_wea_delay,
        addra_out     => AS_L5PHICn2_writeaddr_delay,
        dina_out      => AS_L5PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L5PHICn2_start
      );

    AS_L5PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIDn2_wea_delay,
        addra     => AS_L5PHIDn2_writeaddr_delay,
        dina      => AS_L5PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIDn2_V_readaddr,
        doutb     => AS_L5PHIDn2_V_dout,
        sync_nent => AS_L5PHIDn2_start,
        nent_o    => open
      );

    AS_L5PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIDn2_wea,
        addra     => AS_L5PHIDn2_writeaddr,
        dina      => AS_L5PHIDn2_din,
        wea_out       => AS_L5PHIDn2_wea_delay,
        addra_out     => AS_L5PHIDn2_writeaddr_delay,
        dina_out      => AS_L5PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L5PHIDn2_start
      );

    AS_L6PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIAn2_wea_delay,
        addra     => AS_L6PHIAn2_writeaddr_delay,
        dina      => AS_L6PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIAn2_V_readaddr,
        doutb     => AS_L6PHIAn2_V_dout,
        sync_nent => AS_L6PHIAn2_start,
        nent_o    => open
      );

    AS_L6PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIAn2_wea,
        addra     => AS_L6PHIAn2_writeaddr,
        dina      => AS_L6PHIAn2_din,
        wea_out       => AS_L6PHIAn2_wea_delay,
        addra_out     => AS_L6PHIAn2_writeaddr_delay,
        dina_out      => AS_L6PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_L6PHIAn2_start
      );

    AS_L6PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIBn2_wea_delay,
        addra     => AS_L6PHIBn2_writeaddr_delay,
        dina      => AS_L6PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIBn2_V_readaddr,
        doutb     => AS_L6PHIBn2_V_dout,
        sync_nent => AS_L6PHIBn2_start,
        nent_o    => open
      );

    AS_L6PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIBn2_wea,
        addra     => AS_L6PHIBn2_writeaddr,
        dina      => AS_L6PHIBn2_din,
        wea_out       => AS_L6PHIBn2_wea_delay,
        addra_out     => AS_L6PHIBn2_writeaddr_delay,
        dina_out      => AS_L6PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_L6PHIBn2_start
      );

    AS_L6PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHICn2_wea_delay,
        addra     => AS_L6PHICn2_writeaddr_delay,
        dina      => AS_L6PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHICn2_V_readaddr,
        doutb     => AS_L6PHICn2_V_dout,
        sync_nent => AS_L6PHICn2_start,
        nent_o    => open
      );

    AS_L6PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHICn2_wea,
        addra     => AS_L6PHICn2_writeaddr,
        dina      => AS_L6PHICn2_din,
        wea_out       => AS_L6PHICn2_wea_delay,
        addra_out     => AS_L6PHICn2_writeaddr_delay,
        dina_out      => AS_L6PHICn2_din_delay,
        done       => PC_done,
        start      => AS_L6PHICn2_start
      );

    AS_L6PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIDn2_wea_delay,
        addra     => AS_L6PHIDn2_writeaddr_delay,
        dina      => AS_L6PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIDn2_V_readaddr,
        doutb     => AS_L6PHIDn2_V_dout,
        sync_nent => AS_L6PHIDn2_start,
        nent_o    => open
      );

    AS_L6PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIDn2_wea,
        addra     => AS_L6PHIDn2_writeaddr,
        dina      => AS_L6PHIDn2_din,
        wea_out       => AS_L6PHIDn2_wea_delay,
        addra_out     => AS_L6PHIDn2_writeaddr_delay,
        dina_out      => AS_L6PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_L6PHIDn2_start
      );

    AS_D1PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIAn2_wea_delay,
        addra     => AS_D1PHIAn2_writeaddr_delay,
        dina      => AS_D1PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIAn2_V_readaddr,
        doutb     => AS_D1PHIAn2_V_dout,
        sync_nent => AS_D1PHIAn2_start,
        nent_o    => open
      );

    AS_D1PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIAn2_wea,
        addra     => AS_D1PHIAn2_writeaddr,
        dina      => AS_D1PHIAn2_din,
        wea_out       => AS_D1PHIAn2_wea_delay,
        addra_out     => AS_D1PHIAn2_writeaddr_delay,
        dina_out      => AS_D1PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_D1PHIAn2_start
      );

    AS_D1PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIBn2_wea_delay,
        addra     => AS_D1PHIBn2_writeaddr_delay,
        dina      => AS_D1PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIBn2_V_readaddr,
        doutb     => AS_D1PHIBn2_V_dout,
        sync_nent => AS_D1PHIBn2_start,
        nent_o    => open
      );

    AS_D1PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIBn2_wea,
        addra     => AS_D1PHIBn2_writeaddr,
        dina      => AS_D1PHIBn2_din,
        wea_out       => AS_D1PHIBn2_wea_delay,
        addra_out     => AS_D1PHIBn2_writeaddr_delay,
        dina_out      => AS_D1PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_D1PHIBn2_start
      );

    AS_D1PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHICn2_wea_delay,
        addra     => AS_D1PHICn2_writeaddr_delay,
        dina      => AS_D1PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHICn2_V_readaddr,
        doutb     => AS_D1PHICn2_V_dout,
        sync_nent => AS_D1PHICn2_start,
        nent_o    => open
      );

    AS_D1PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHICn2_wea,
        addra     => AS_D1PHICn2_writeaddr,
        dina      => AS_D1PHICn2_din,
        wea_out       => AS_D1PHICn2_wea_delay,
        addra_out     => AS_D1PHICn2_writeaddr_delay,
        dina_out      => AS_D1PHICn2_din_delay,
        done       => PC_done,
        start      => AS_D1PHICn2_start
      );

    AS_D1PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIDn2_wea_delay,
        addra     => AS_D1PHIDn2_writeaddr_delay,
        dina      => AS_D1PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIDn2_V_readaddr,
        doutb     => AS_D1PHIDn2_V_dout,
        sync_nent => AS_D1PHIDn2_start,
        nent_o    => open
      );

    AS_D1PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIDn2_wea,
        addra     => AS_D1PHIDn2_writeaddr,
        dina      => AS_D1PHIDn2_din,
        wea_out       => AS_D1PHIDn2_wea_delay,
        addra_out     => AS_D1PHIDn2_writeaddr_delay,
        dina_out      => AS_D1PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_D1PHIDn2_start
      );

    AS_D2PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIAn2_wea_delay,
        addra     => AS_D2PHIAn2_writeaddr_delay,
        dina      => AS_D2PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIAn2_V_readaddr,
        doutb     => AS_D2PHIAn2_V_dout,
        sync_nent => AS_D2PHIAn2_start,
        nent_o    => open
      );

    AS_D2PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIAn2_wea,
        addra     => AS_D2PHIAn2_writeaddr,
        dina      => AS_D2PHIAn2_din,
        wea_out       => AS_D2PHIAn2_wea_delay,
        addra_out     => AS_D2PHIAn2_writeaddr_delay,
        dina_out      => AS_D2PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_D2PHIAn2_start
      );

    AS_D2PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIBn2_wea_delay,
        addra     => AS_D2PHIBn2_writeaddr_delay,
        dina      => AS_D2PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIBn2_V_readaddr,
        doutb     => AS_D2PHIBn2_V_dout,
        sync_nent => AS_D2PHIBn2_start,
        nent_o    => open
      );

    AS_D2PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIBn2_wea,
        addra     => AS_D2PHIBn2_writeaddr,
        dina      => AS_D2PHIBn2_din,
        wea_out       => AS_D2PHIBn2_wea_delay,
        addra_out     => AS_D2PHIBn2_writeaddr_delay,
        dina_out      => AS_D2PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_D2PHIBn2_start
      );

    AS_D2PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHICn2_wea_delay,
        addra     => AS_D2PHICn2_writeaddr_delay,
        dina      => AS_D2PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHICn2_V_readaddr,
        doutb     => AS_D2PHICn2_V_dout,
        sync_nent => AS_D2PHICn2_start,
        nent_o    => open
      );

    AS_D2PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHICn2_wea,
        addra     => AS_D2PHICn2_writeaddr,
        dina      => AS_D2PHICn2_din,
        wea_out       => AS_D2PHICn2_wea_delay,
        addra_out     => AS_D2PHICn2_writeaddr_delay,
        dina_out      => AS_D2PHICn2_din_delay,
        done       => PC_done,
        start      => AS_D2PHICn2_start
      );

    AS_D2PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIDn2_wea_delay,
        addra     => AS_D2PHIDn2_writeaddr_delay,
        dina      => AS_D2PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIDn2_V_readaddr,
        doutb     => AS_D2PHIDn2_V_dout,
        sync_nent => AS_D2PHIDn2_start,
        nent_o    => open
      );

    AS_D2PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIDn2_wea,
        addra     => AS_D2PHIDn2_writeaddr,
        dina      => AS_D2PHIDn2_din,
        wea_out       => AS_D2PHIDn2_wea_delay,
        addra_out     => AS_D2PHIDn2_writeaddr_delay,
        dina_out      => AS_D2PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_D2PHIDn2_start
      );

    AS_D3PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIAn2_wea_delay,
        addra     => AS_D3PHIAn2_writeaddr_delay,
        dina      => AS_D3PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIAn2_V_readaddr,
        doutb     => AS_D3PHIAn2_V_dout,
        sync_nent => AS_D3PHIAn2_start,
        nent_o    => open
      );

    AS_D3PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIAn2_wea,
        addra     => AS_D3PHIAn2_writeaddr,
        dina      => AS_D3PHIAn2_din,
        wea_out       => AS_D3PHIAn2_wea_delay,
        addra_out     => AS_D3PHIAn2_writeaddr_delay,
        dina_out      => AS_D3PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_D3PHIAn2_start
      );

    AS_D3PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIBn2_wea_delay,
        addra     => AS_D3PHIBn2_writeaddr_delay,
        dina      => AS_D3PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIBn2_V_readaddr,
        doutb     => AS_D3PHIBn2_V_dout,
        sync_nent => AS_D3PHIBn2_start,
        nent_o    => open
      );

    AS_D3PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIBn2_wea,
        addra     => AS_D3PHIBn2_writeaddr,
        dina      => AS_D3PHIBn2_din,
        wea_out       => AS_D3PHIBn2_wea_delay,
        addra_out     => AS_D3PHIBn2_writeaddr_delay,
        dina_out      => AS_D3PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_D3PHIBn2_start
      );

    AS_D3PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHICn2_wea_delay,
        addra     => AS_D3PHICn2_writeaddr_delay,
        dina      => AS_D3PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHICn2_V_readaddr,
        doutb     => AS_D3PHICn2_V_dout,
        sync_nent => AS_D3PHICn2_start,
        nent_o    => open
      );

    AS_D3PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHICn2_wea,
        addra     => AS_D3PHICn2_writeaddr,
        dina      => AS_D3PHICn2_din,
        wea_out       => AS_D3PHICn2_wea_delay,
        addra_out     => AS_D3PHICn2_writeaddr_delay,
        dina_out      => AS_D3PHICn2_din_delay,
        done       => PC_done,
        start      => AS_D3PHICn2_start
      );

    AS_D3PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIDn2_wea_delay,
        addra     => AS_D3PHIDn2_writeaddr_delay,
        dina      => AS_D3PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIDn2_V_readaddr,
        doutb     => AS_D3PHIDn2_V_dout,
        sync_nent => AS_D3PHIDn2_start,
        nent_o    => open
      );

    AS_D3PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIDn2_wea,
        addra     => AS_D3PHIDn2_writeaddr,
        dina      => AS_D3PHIDn2_din,
        wea_out       => AS_D3PHIDn2_wea_delay,
        addra_out     => AS_D3PHIDn2_writeaddr_delay,
        dina_out      => AS_D3PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_D3PHIDn2_start
      );

    AS_D4PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIAn2_wea_delay,
        addra     => AS_D4PHIAn2_writeaddr_delay,
        dina      => AS_D4PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIAn2_V_readaddr,
        doutb     => AS_D4PHIAn2_V_dout,
        sync_nent => AS_D4PHIAn2_start,
        nent_o    => open
      );

    AS_D4PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIAn2_wea,
        addra     => AS_D4PHIAn2_writeaddr,
        dina      => AS_D4PHIAn2_din,
        wea_out       => AS_D4PHIAn2_wea_delay,
        addra_out     => AS_D4PHIAn2_writeaddr_delay,
        dina_out      => AS_D4PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_D4PHIAn2_start
      );

    AS_D4PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIBn2_wea_delay,
        addra     => AS_D4PHIBn2_writeaddr_delay,
        dina      => AS_D4PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIBn2_V_readaddr,
        doutb     => AS_D4PHIBn2_V_dout,
        sync_nent => AS_D4PHIBn2_start,
        nent_o    => open
      );

    AS_D4PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIBn2_wea,
        addra     => AS_D4PHIBn2_writeaddr,
        dina      => AS_D4PHIBn2_din,
        wea_out       => AS_D4PHIBn2_wea_delay,
        addra_out     => AS_D4PHIBn2_writeaddr_delay,
        dina_out      => AS_D4PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_D4PHIBn2_start
      );

    AS_D4PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHICn2_wea_delay,
        addra     => AS_D4PHICn2_writeaddr_delay,
        dina      => AS_D4PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHICn2_V_readaddr,
        doutb     => AS_D4PHICn2_V_dout,
        sync_nent => AS_D4PHICn2_start,
        nent_o    => open
      );

    AS_D4PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHICn2_wea,
        addra     => AS_D4PHICn2_writeaddr,
        dina      => AS_D4PHICn2_din,
        wea_out       => AS_D4PHICn2_wea_delay,
        addra_out     => AS_D4PHICn2_writeaddr_delay,
        dina_out      => AS_D4PHICn2_din_delay,
        done       => PC_done,
        start      => AS_D4PHICn2_start
      );

    AS_D4PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIDn2_wea_delay,
        addra     => AS_D4PHIDn2_writeaddr_delay,
        dina      => AS_D4PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIDn2_V_readaddr,
        doutb     => AS_D4PHIDn2_V_dout,
        sync_nent => AS_D4PHIDn2_start,
        nent_o    => open
      );

    AS_D4PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIDn2_wea,
        addra     => AS_D4PHIDn2_writeaddr,
        dina      => AS_D4PHIDn2_din,
        wea_out       => AS_D4PHIDn2_wea_delay,
        addra_out     => AS_D4PHIDn2_writeaddr_delay,
        dina_out      => AS_D4PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_D4PHIDn2_start
      );

    AS_D5PHIAn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIAn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIAn2_wea_delay,
        addra     => AS_D5PHIAn2_writeaddr_delay,
        dina      => AS_D5PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIAn2_V_readaddr,
        doutb     => AS_D5PHIAn2_V_dout,
        sync_nent => AS_D5PHIAn2_start,
        nent_o    => open
      );

    AS_D5PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIAn2_wea,
        addra     => AS_D5PHIAn2_writeaddr,
        dina      => AS_D5PHIAn2_din,
        wea_out       => AS_D5PHIAn2_wea_delay,
        addra_out     => AS_D5PHIAn2_writeaddr_delay,
        dina_out      => AS_D5PHIAn2_din_delay,
        done       => PC_done,
        start      => AS_D5PHIAn2_start
      );

    AS_D5PHIBn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIBn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIBn2_wea_delay,
        addra     => AS_D5PHIBn2_writeaddr_delay,
        dina      => AS_D5PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIBn2_V_readaddr,
        doutb     => AS_D5PHIBn2_V_dout,
        sync_nent => AS_D5PHIBn2_start,
        nent_o    => open
      );

    AS_D5PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIBn2_wea,
        addra     => AS_D5PHIBn2_writeaddr,
        dina      => AS_D5PHIBn2_din,
        wea_out       => AS_D5PHIBn2_wea_delay,
        addra_out     => AS_D5PHIBn2_writeaddr_delay,
        dina_out      => AS_D5PHIBn2_din_delay,
        done       => PC_done,
        start      => AS_D5PHIBn2_start
      );

    AS_D5PHICn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHICn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHICn2_wea_delay,
        addra     => AS_D5PHICn2_writeaddr_delay,
        dina      => AS_D5PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHICn2_V_readaddr,
        doutb     => AS_D5PHICn2_V_dout,
        sync_nent => AS_D5PHICn2_start,
        nent_o    => open
      );

    AS_D5PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHICn2_wea,
        addra     => AS_D5PHICn2_writeaddr,
        dina      => AS_D5PHICn2_din,
        wea_out       => AS_D5PHICn2_wea_delay,
        addra_out     => AS_D5PHICn2_writeaddr_delay,
        dina_out      => AS_D5PHICn2_din_delay,
        done       => PC_done,
        start      => AS_D5PHICn2_start
      );

    AS_D5PHIDn2 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIDn2"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIDn2_wea_delay,
        addra     => AS_D5PHIDn2_writeaddr_delay,
        dina      => AS_D5PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIDn2_V_readaddr,
        doutb     => AS_D5PHIDn2_V_dout,
        sync_nent => AS_D5PHIDn2_start,
        nent_o    => open
      );

    AS_D5PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIDn2_wea,
        addra     => AS_D5PHIDn2_writeaddr,
        dina      => AS_D5PHIDn2_din,
        wea_out       => AS_D5PHIDn2_wea_delay,
        addra_out     => AS_D5PHIDn2_writeaddr_delay,
        dina_out      => AS_D5PHIDn2_din_delay,
        done       => PC_done,
        start      => AS_D5PHIDn2_start
      );

    VMSME_L1PHIAn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIAn2_V_datatmp,
        dataout0 => VMSME_L1PHIAn2_AV_dout(0),
        dataout1 => VMSME_L1PHIAn2_AV_dout(1),
        dataout2 => VMSME_L1PHIAn2_AV_dout(2),
        dataout3 => VMSME_L1PHIAn2_AV_dout(3)
      );

    VMSME_L1PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIAn2_wea_delay,
        addra     => VMSME_L1PHIAn2_writeaddr_delay,
        dina      => VMSME_L1PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIAn2_AV_readaddr(3),VMSME_L1PHIAn2_AV_readaddr(2),VMSME_L1PHIAn2_AV_readaddr(1),VMSME_L1PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIAn2_V_datatmp,
        enb_nent  => VMSME_L1PHIAn2_enb_nent,
        addr_nent  => VMSME_L1PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIAn2_V_binmaskb
      );

    VMSME_L1PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIAn2_wea,
        addra     => VMSME_L1PHIAn2_writeaddr,
        dina      => VMSME_L1PHIAn2_din,
        wea_out       => VMSME_L1PHIAn2_wea_delay,
        addra_out     => VMSME_L1PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIAn2_start
      );

    VMSME_L1PHIBn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIBn2_V_datatmp,
        dataout0 => VMSME_L1PHIBn2_AV_dout(0),
        dataout1 => VMSME_L1PHIBn2_AV_dout(1),
        dataout2 => VMSME_L1PHIBn2_AV_dout(2),
        dataout3 => VMSME_L1PHIBn2_AV_dout(3)
      );

    VMSME_L1PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIBn2_wea_delay,
        addra     => VMSME_L1PHIBn2_writeaddr_delay,
        dina      => VMSME_L1PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIBn2_AV_readaddr(3),VMSME_L1PHIBn2_AV_readaddr(2),VMSME_L1PHIBn2_AV_readaddr(1),VMSME_L1PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIBn2_V_datatmp,
        enb_nent  => VMSME_L1PHIBn2_enb_nent,
        addr_nent  => VMSME_L1PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIBn2_V_binmaskb
      );

    VMSME_L1PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIBn2_wea,
        addra     => VMSME_L1PHIBn2_writeaddr,
        dina      => VMSME_L1PHIBn2_din,
        wea_out       => VMSME_L1PHIBn2_wea_delay,
        addra_out     => VMSME_L1PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIBn2_start
      );

    VMSME_L1PHICn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHICn2_V_datatmp,
        dataout0 => VMSME_L1PHICn2_AV_dout(0),
        dataout1 => VMSME_L1PHICn2_AV_dout(1),
        dataout2 => VMSME_L1PHICn2_AV_dout(2),
        dataout3 => VMSME_L1PHICn2_AV_dout(3)
      );

    VMSME_L1PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHICn2_wea_delay,
        addra     => VMSME_L1PHICn2_writeaddr_delay,
        dina      => VMSME_L1PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHICn2_AV_readaddr(3),VMSME_L1PHICn2_AV_readaddr(2),VMSME_L1PHICn2_AV_readaddr(1),VMSME_L1PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHICn2_V_datatmp,
        enb_nent  => VMSME_L1PHICn2_enb_nent,
        addr_nent  => VMSME_L1PHICn2_V_addr_nent,
        dout_nent  => VMSME_L1PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHICn2_V_binmaskb
      );

    VMSME_L1PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHICn2_wea,
        addra     => VMSME_L1PHICn2_writeaddr,
        dina      => VMSME_L1PHICn2_din,
        wea_out       => VMSME_L1PHICn2_wea_delay,
        addra_out     => VMSME_L1PHICn2_writeaddr_delay,
        dina_out      => VMSME_L1PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHICn2_start
      );

    VMSME_L1PHIDn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIDn2_V_datatmp,
        dataout0 => VMSME_L1PHIDn2_AV_dout(0),
        dataout1 => VMSME_L1PHIDn2_AV_dout(1),
        dataout2 => VMSME_L1PHIDn2_AV_dout(2),
        dataout3 => VMSME_L1PHIDn2_AV_dout(3)
      );

    VMSME_L1PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIDn2_wea_delay,
        addra     => VMSME_L1PHIDn2_writeaddr_delay,
        dina      => VMSME_L1PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIDn2_AV_readaddr(3),VMSME_L1PHIDn2_AV_readaddr(2),VMSME_L1PHIDn2_AV_readaddr(1),VMSME_L1PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIDn2_V_datatmp,
        enb_nent  => VMSME_L1PHIDn2_enb_nent,
        addr_nent  => VMSME_L1PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIDn2_V_binmaskb
      );

    VMSME_L1PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIDn2_wea,
        addra     => VMSME_L1PHIDn2_writeaddr,
        dina      => VMSME_L1PHIDn2_din,
        wea_out       => VMSME_L1PHIDn2_wea_delay,
        addra_out     => VMSME_L1PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIDn2_start
      );

    VMSME_L1PHIEn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIEn2_V_datatmp,
        dataout0 => VMSME_L1PHIEn2_AV_dout(0),
        dataout1 => VMSME_L1PHIEn2_AV_dout(1),
        dataout2 => VMSME_L1PHIEn2_AV_dout(2),
        dataout3 => VMSME_L1PHIEn2_AV_dout(3)
      );

    VMSME_L1PHIEn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIEn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIEn2_wea_delay,
        addra     => VMSME_L1PHIEn2_writeaddr_delay,
        dina      => VMSME_L1PHIEn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIEn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIEn2_AV_readaddr(3),VMSME_L1PHIEn2_AV_readaddr(2),VMSME_L1PHIEn2_AV_readaddr(1),VMSME_L1PHIEn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIEn2_V_datatmp,
        enb_nent  => VMSME_L1PHIEn2_enb_nent,
        addr_nent  => VMSME_L1PHIEn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIEn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIEn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIEn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIEn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIEn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIEn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIEn2_V_binmaskb
      );

    VMSME_L1PHIEn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIEn2_wea,
        addra     => VMSME_L1PHIEn2_writeaddr,
        dina      => VMSME_L1PHIEn2_din,
        wea_out       => VMSME_L1PHIEn2_wea_delay,
        addra_out     => VMSME_L1PHIEn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIEn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIEn2_start
      );

    VMSME_L1PHIFn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIFn2_V_datatmp,
        dataout0 => VMSME_L1PHIFn2_AV_dout(0),
        dataout1 => VMSME_L1PHIFn2_AV_dout(1),
        dataout2 => VMSME_L1PHIFn2_AV_dout(2),
        dataout3 => VMSME_L1PHIFn2_AV_dout(3)
      );

    VMSME_L1PHIFn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIFn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIFn2_wea_delay,
        addra     => VMSME_L1PHIFn2_writeaddr_delay,
        dina      => VMSME_L1PHIFn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIFn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIFn2_AV_readaddr(3),VMSME_L1PHIFn2_AV_readaddr(2),VMSME_L1PHIFn2_AV_readaddr(1),VMSME_L1PHIFn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIFn2_V_datatmp,
        enb_nent  => VMSME_L1PHIFn2_enb_nent,
        addr_nent  => VMSME_L1PHIFn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIFn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIFn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIFn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIFn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIFn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIFn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIFn2_V_binmaskb
      );

    VMSME_L1PHIFn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIFn2_wea,
        addra     => VMSME_L1PHIFn2_writeaddr,
        dina      => VMSME_L1PHIFn2_din,
        wea_out       => VMSME_L1PHIFn2_wea_delay,
        addra_out     => VMSME_L1PHIFn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIFn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIFn2_start
      );

    VMSME_L1PHIGn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIGn2_V_datatmp,
        dataout0 => VMSME_L1PHIGn2_AV_dout(0),
        dataout1 => VMSME_L1PHIGn2_AV_dout(1),
        dataout2 => VMSME_L1PHIGn2_AV_dout(2),
        dataout3 => VMSME_L1PHIGn2_AV_dout(3)
      );

    VMSME_L1PHIGn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIGn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIGn2_wea_delay,
        addra     => VMSME_L1PHIGn2_writeaddr_delay,
        dina      => VMSME_L1PHIGn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIGn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIGn2_AV_readaddr(3),VMSME_L1PHIGn2_AV_readaddr(2),VMSME_L1PHIGn2_AV_readaddr(1),VMSME_L1PHIGn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIGn2_V_datatmp,
        enb_nent  => VMSME_L1PHIGn2_enb_nent,
        addr_nent  => VMSME_L1PHIGn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIGn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIGn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIGn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIGn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIGn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIGn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIGn2_V_binmaskb
      );

    VMSME_L1PHIGn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIGn2_wea,
        addra     => VMSME_L1PHIGn2_writeaddr,
        dina      => VMSME_L1PHIGn2_din,
        wea_out       => VMSME_L1PHIGn2_wea_delay,
        addra_out     => VMSME_L1PHIGn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIGn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIGn2_start
      );

    VMSME_L1PHIHn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L1PHIHn2_V_datatmp,
        dataout0 => VMSME_L1PHIHn2_AV_dout(0),
        dataout1 => VMSME_L1PHIHn2_AV_dout(1),
        dataout2 => VMSME_L1PHIHn2_AV_dout(2),
        dataout3 => VMSME_L1PHIHn2_AV_dout(3)
      );

    VMSME_L1PHIHn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L1PHIHn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L1PHIHn2_wea_delay,
        addra     => VMSME_L1PHIHn2_writeaddr_delay,
        dina      => VMSME_L1PHIHn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L1PHIHn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L1PHIHn2_AV_readaddr(3),VMSME_L1PHIHn2_AV_readaddr(2),VMSME_L1PHIHn2_AV_readaddr(1),VMSME_L1PHIHn2_AV_readaddr(0)),
        doutb     => VMSME_L1PHIHn2_V_datatmp,
        enb_nent  => VMSME_L1PHIHn2_enb_nent,
        addr_nent  => VMSME_L1PHIHn2_V_addr_nent,
        dout_nent  => VMSME_L1PHIHn2_AV_dout_nent,
        enb_binmaska  => VMSME_L1PHIHn2_enb_binmaska,
        addr_binmaska  => VMSME_L1PHIHn2_V_addr_binmaska,
        binmaska_o  => VMSME_L1PHIHn2_V_binmaska,
        enb_binmaskb  => VMSME_L1PHIHn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L1PHIHn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L1PHIHn2_V_binmaskb
      );

    VMSME_L1PHIHn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L1PHIHn2_wea,
        addra     => VMSME_L1PHIHn2_writeaddr,
        dina      => VMSME_L1PHIHn2_din,
        wea_out       => VMSME_L1PHIHn2_wea_delay,
        addra_out     => VMSME_L1PHIHn2_writeaddr_delay,
        dina_out      => VMSME_L1PHIHn2_din_delay,
        done       => PC_done,
        start      => VMSME_L1PHIHn2_start
      );

    VMSME_L2PHIAn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L2PHIAn2_V_datatmp,
        dataout0 => VMSME_L2PHIAn2_AV_dout(0),
        dataout1 => VMSME_L2PHIAn2_AV_dout(1),
        dataout2 => VMSME_L2PHIAn2_AV_dout(2),
        dataout3 => VMSME_L2PHIAn2_AV_dout(3)
      );

    VMSME_L2PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L2PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L2PHIAn2_wea_delay,
        addra     => VMSME_L2PHIAn2_writeaddr_delay,
        dina      => VMSME_L2PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L2PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L2PHIAn2_AV_readaddr(3),VMSME_L2PHIAn2_AV_readaddr(2),VMSME_L2PHIAn2_AV_readaddr(1),VMSME_L2PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L2PHIAn2_V_datatmp,
        enb_nent  => VMSME_L2PHIAn2_enb_nent,
        addr_nent  => VMSME_L2PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L2PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L2PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L2PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L2PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L2PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L2PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L2PHIAn2_V_binmaskb
      );

    VMSME_L2PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L2PHIAn2_wea,
        addra     => VMSME_L2PHIAn2_writeaddr,
        dina      => VMSME_L2PHIAn2_din,
        wea_out       => VMSME_L2PHIAn2_wea_delay,
        addra_out     => VMSME_L2PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L2PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L2PHIAn2_start
      );

    VMSME_L2PHIBn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L2PHIBn2_V_datatmp,
        dataout0 => VMSME_L2PHIBn2_AV_dout(0),
        dataout1 => VMSME_L2PHIBn2_AV_dout(1),
        dataout2 => VMSME_L2PHIBn2_AV_dout(2),
        dataout3 => VMSME_L2PHIBn2_AV_dout(3)
      );

    VMSME_L2PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L2PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L2PHIBn2_wea_delay,
        addra     => VMSME_L2PHIBn2_writeaddr_delay,
        dina      => VMSME_L2PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L2PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L2PHIBn2_AV_readaddr(3),VMSME_L2PHIBn2_AV_readaddr(2),VMSME_L2PHIBn2_AV_readaddr(1),VMSME_L2PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L2PHIBn2_V_datatmp,
        enb_nent  => VMSME_L2PHIBn2_enb_nent,
        addr_nent  => VMSME_L2PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L2PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L2PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L2PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L2PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L2PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L2PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L2PHIBn2_V_binmaskb
      );

    VMSME_L2PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L2PHIBn2_wea,
        addra     => VMSME_L2PHIBn2_writeaddr,
        dina      => VMSME_L2PHIBn2_din,
        wea_out       => VMSME_L2PHIBn2_wea_delay,
        addra_out     => VMSME_L2PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L2PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L2PHIBn2_start
      );

    VMSME_L2PHICn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L2PHICn2_V_datatmp,
        dataout0 => VMSME_L2PHICn2_AV_dout(0),
        dataout1 => VMSME_L2PHICn2_AV_dout(1),
        dataout2 => VMSME_L2PHICn2_AV_dout(2),
        dataout3 => VMSME_L2PHICn2_AV_dout(3)
      );

    VMSME_L2PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L2PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L2PHICn2_wea_delay,
        addra     => VMSME_L2PHICn2_writeaddr_delay,
        dina      => VMSME_L2PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L2PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L2PHICn2_AV_readaddr(3),VMSME_L2PHICn2_AV_readaddr(2),VMSME_L2PHICn2_AV_readaddr(1),VMSME_L2PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L2PHICn2_V_datatmp,
        enb_nent  => VMSME_L2PHICn2_enb_nent,
        addr_nent  => VMSME_L2PHICn2_V_addr_nent,
        dout_nent  => VMSME_L2PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L2PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L2PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L2PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L2PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L2PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L2PHICn2_V_binmaskb
      );

    VMSME_L2PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L2PHICn2_wea,
        addra     => VMSME_L2PHICn2_writeaddr,
        dina      => VMSME_L2PHICn2_din,
        wea_out       => VMSME_L2PHICn2_wea_delay,
        addra_out     => VMSME_L2PHICn2_writeaddr_delay,
        dina_out      => VMSME_L2PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L2PHICn2_start
      );

    VMSME_L2PHIDn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L2PHIDn2_V_datatmp,
        dataout0 => VMSME_L2PHIDn2_AV_dout(0),
        dataout1 => VMSME_L2PHIDn2_AV_dout(1),
        dataout2 => VMSME_L2PHIDn2_AV_dout(2),
        dataout3 => VMSME_L2PHIDn2_AV_dout(3)
      );

    VMSME_L2PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L2PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L2PHIDn2_wea_delay,
        addra     => VMSME_L2PHIDn2_writeaddr_delay,
        dina      => VMSME_L2PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L2PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L2PHIDn2_AV_readaddr(3),VMSME_L2PHIDn2_AV_readaddr(2),VMSME_L2PHIDn2_AV_readaddr(1),VMSME_L2PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L2PHIDn2_V_datatmp,
        enb_nent  => VMSME_L2PHIDn2_enb_nent,
        addr_nent  => VMSME_L2PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L2PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L2PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L2PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L2PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L2PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L2PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L2PHIDn2_V_binmaskb
      );

    VMSME_L2PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L2PHIDn2_wea,
        addra     => VMSME_L2PHIDn2_writeaddr,
        dina      => VMSME_L2PHIDn2_din,
        wea_out       => VMSME_L2PHIDn2_wea_delay,
        addra_out     => VMSME_L2PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L2PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L2PHIDn2_start
      );

    VMSME_L3PHIAn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L3PHIAn2_V_datatmp,
        dataout0 => VMSME_L3PHIAn2_AV_dout(0),
        dataout1 => VMSME_L3PHIAn2_AV_dout(1),
        dataout2 => VMSME_L3PHIAn2_AV_dout(2),
        dataout3 => VMSME_L3PHIAn2_AV_dout(3)
      );

    VMSME_L3PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L3PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L3PHIAn2_wea_delay,
        addra     => VMSME_L3PHIAn2_writeaddr_delay,
        dina      => VMSME_L3PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L3PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L3PHIAn2_AV_readaddr(3),VMSME_L3PHIAn2_AV_readaddr(2),VMSME_L3PHIAn2_AV_readaddr(1),VMSME_L3PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L3PHIAn2_V_datatmp,
        enb_nent  => VMSME_L3PHIAn2_enb_nent,
        addr_nent  => VMSME_L3PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L3PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L3PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L3PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L3PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L3PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L3PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L3PHIAn2_V_binmaskb
      );

    VMSME_L3PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L3PHIAn2_wea,
        addra     => VMSME_L3PHIAn2_writeaddr,
        dina      => VMSME_L3PHIAn2_din,
        wea_out       => VMSME_L3PHIAn2_wea_delay,
        addra_out     => VMSME_L3PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L3PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L3PHIAn2_start
      );

    VMSME_L3PHIBn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L3PHIBn2_V_datatmp,
        dataout0 => VMSME_L3PHIBn2_AV_dout(0),
        dataout1 => VMSME_L3PHIBn2_AV_dout(1),
        dataout2 => VMSME_L3PHIBn2_AV_dout(2),
        dataout3 => VMSME_L3PHIBn2_AV_dout(3)
      );

    VMSME_L3PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L3PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L3PHIBn2_wea_delay,
        addra     => VMSME_L3PHIBn2_writeaddr_delay,
        dina      => VMSME_L3PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L3PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L3PHIBn2_AV_readaddr(3),VMSME_L3PHIBn2_AV_readaddr(2),VMSME_L3PHIBn2_AV_readaddr(1),VMSME_L3PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L3PHIBn2_V_datatmp,
        enb_nent  => VMSME_L3PHIBn2_enb_nent,
        addr_nent  => VMSME_L3PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L3PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L3PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L3PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L3PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L3PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L3PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L3PHIBn2_V_binmaskb
      );

    VMSME_L3PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L3PHIBn2_wea,
        addra     => VMSME_L3PHIBn2_writeaddr,
        dina      => VMSME_L3PHIBn2_din,
        wea_out       => VMSME_L3PHIBn2_wea_delay,
        addra_out     => VMSME_L3PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L3PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L3PHIBn2_start
      );

    VMSME_L3PHICn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L3PHICn2_V_datatmp,
        dataout0 => VMSME_L3PHICn2_AV_dout(0),
        dataout1 => VMSME_L3PHICn2_AV_dout(1),
        dataout2 => VMSME_L3PHICn2_AV_dout(2),
        dataout3 => VMSME_L3PHICn2_AV_dout(3)
      );

    VMSME_L3PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L3PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L3PHICn2_wea_delay,
        addra     => VMSME_L3PHICn2_writeaddr_delay,
        dina      => VMSME_L3PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L3PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L3PHICn2_AV_readaddr(3),VMSME_L3PHICn2_AV_readaddr(2),VMSME_L3PHICn2_AV_readaddr(1),VMSME_L3PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L3PHICn2_V_datatmp,
        enb_nent  => VMSME_L3PHICn2_enb_nent,
        addr_nent  => VMSME_L3PHICn2_V_addr_nent,
        dout_nent  => VMSME_L3PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L3PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L3PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L3PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L3PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L3PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L3PHICn2_V_binmaskb
      );

    VMSME_L3PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L3PHICn2_wea,
        addra     => VMSME_L3PHICn2_writeaddr,
        dina      => VMSME_L3PHICn2_din,
        wea_out       => VMSME_L3PHICn2_wea_delay,
        addra_out     => VMSME_L3PHICn2_writeaddr_delay,
        dina_out      => VMSME_L3PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L3PHICn2_start
      );

    VMSME_L3PHIDn2_dataformat : entity work.vmstub16dout4
      port map (
        datain => VMSME_L3PHIDn2_V_datatmp,
        dataout0 => VMSME_L3PHIDn2_AV_dout(0),
        dataout1 => VMSME_L3PHIDn2_AV_dout(1),
        dataout2 => VMSME_L3PHIDn2_AV_dout(2),
        dataout3 => VMSME_L3PHIDn2_AV_dout(3)
      );

    VMSME_L3PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L3PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L3PHIDn2_wea_delay,
        addra     => VMSME_L3PHIDn2_writeaddr_delay,
        dina      => VMSME_L3PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L3PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L3PHIDn2_AV_readaddr(3),VMSME_L3PHIDn2_AV_readaddr(2),VMSME_L3PHIDn2_AV_readaddr(1),VMSME_L3PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L3PHIDn2_V_datatmp,
        enb_nent  => VMSME_L3PHIDn2_enb_nent,
        addr_nent  => VMSME_L3PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L3PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L3PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L3PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L3PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L3PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L3PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L3PHIDn2_V_binmaskb
      );

    VMSME_L3PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSME_L3PHIDn2_wea,
        addra     => VMSME_L3PHIDn2_writeaddr,
        dina      => VMSME_L3PHIDn2_din,
        wea_out       => VMSME_L3PHIDn2_wea_delay,
        addra_out     => VMSME_L3PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L3PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L3PHIDn2_start
      );

    VMSME_L4PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L4PHIAn2_V_datatmp,
        dataout0 => VMSME_L4PHIAn2_AV_dout(0),
        dataout1 => VMSME_L4PHIAn2_AV_dout(1),
        dataout2 => VMSME_L4PHIAn2_AV_dout(2),
        dataout3 => VMSME_L4PHIAn2_AV_dout(3)
      );

    VMSME_L4PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L4PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L4PHIAn2_wea_delay,
        addra     => VMSME_L4PHIAn2_writeaddr_delay,
        dina      => VMSME_L4PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L4PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L4PHIAn2_AV_readaddr(3),VMSME_L4PHIAn2_AV_readaddr(2),VMSME_L4PHIAn2_AV_readaddr(1),VMSME_L4PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L4PHIAn2_V_datatmp,
        enb_nent  => VMSME_L4PHIAn2_enb_nent,
        addr_nent  => VMSME_L4PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L4PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L4PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L4PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L4PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L4PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L4PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L4PHIAn2_V_binmaskb
      );

    VMSME_L4PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L4PHIAn2_wea,
        addra     => VMSME_L4PHIAn2_writeaddr,
        dina      => VMSME_L4PHIAn2_din,
        wea_out       => VMSME_L4PHIAn2_wea_delay,
        addra_out     => VMSME_L4PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L4PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L4PHIAn2_start
      );

    VMSME_L4PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L4PHIBn2_V_datatmp,
        dataout0 => VMSME_L4PHIBn2_AV_dout(0),
        dataout1 => VMSME_L4PHIBn2_AV_dout(1),
        dataout2 => VMSME_L4PHIBn2_AV_dout(2),
        dataout3 => VMSME_L4PHIBn2_AV_dout(3)
      );

    VMSME_L4PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L4PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L4PHIBn2_wea_delay,
        addra     => VMSME_L4PHIBn2_writeaddr_delay,
        dina      => VMSME_L4PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L4PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L4PHIBn2_AV_readaddr(3),VMSME_L4PHIBn2_AV_readaddr(2),VMSME_L4PHIBn2_AV_readaddr(1),VMSME_L4PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L4PHIBn2_V_datatmp,
        enb_nent  => VMSME_L4PHIBn2_enb_nent,
        addr_nent  => VMSME_L4PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L4PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L4PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L4PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L4PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L4PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L4PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L4PHIBn2_V_binmaskb
      );

    VMSME_L4PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L4PHIBn2_wea,
        addra     => VMSME_L4PHIBn2_writeaddr,
        dina      => VMSME_L4PHIBn2_din,
        wea_out       => VMSME_L4PHIBn2_wea_delay,
        addra_out     => VMSME_L4PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L4PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L4PHIBn2_start
      );

    VMSME_L4PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L4PHICn2_V_datatmp,
        dataout0 => VMSME_L4PHICn2_AV_dout(0),
        dataout1 => VMSME_L4PHICn2_AV_dout(1),
        dataout2 => VMSME_L4PHICn2_AV_dout(2),
        dataout3 => VMSME_L4PHICn2_AV_dout(3)
      );

    VMSME_L4PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L4PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L4PHICn2_wea_delay,
        addra     => VMSME_L4PHICn2_writeaddr_delay,
        dina      => VMSME_L4PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L4PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L4PHICn2_AV_readaddr(3),VMSME_L4PHICn2_AV_readaddr(2),VMSME_L4PHICn2_AV_readaddr(1),VMSME_L4PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L4PHICn2_V_datatmp,
        enb_nent  => VMSME_L4PHICn2_enb_nent,
        addr_nent  => VMSME_L4PHICn2_V_addr_nent,
        dout_nent  => VMSME_L4PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L4PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L4PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L4PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L4PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L4PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L4PHICn2_V_binmaskb
      );

    VMSME_L4PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L4PHICn2_wea,
        addra     => VMSME_L4PHICn2_writeaddr,
        dina      => VMSME_L4PHICn2_din,
        wea_out       => VMSME_L4PHICn2_wea_delay,
        addra_out     => VMSME_L4PHICn2_writeaddr_delay,
        dina_out      => VMSME_L4PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L4PHICn2_start
      );

    VMSME_L4PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L4PHIDn2_V_datatmp,
        dataout0 => VMSME_L4PHIDn2_AV_dout(0),
        dataout1 => VMSME_L4PHIDn2_AV_dout(1),
        dataout2 => VMSME_L4PHIDn2_AV_dout(2),
        dataout3 => VMSME_L4PHIDn2_AV_dout(3)
      );

    VMSME_L4PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L4PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L4PHIDn2_wea_delay,
        addra     => VMSME_L4PHIDn2_writeaddr_delay,
        dina      => VMSME_L4PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L4PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L4PHIDn2_AV_readaddr(3),VMSME_L4PHIDn2_AV_readaddr(2),VMSME_L4PHIDn2_AV_readaddr(1),VMSME_L4PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L4PHIDn2_V_datatmp,
        enb_nent  => VMSME_L4PHIDn2_enb_nent,
        addr_nent  => VMSME_L4PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L4PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L4PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L4PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L4PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L4PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L4PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L4PHIDn2_V_binmaskb
      );

    VMSME_L4PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L4PHIDn2_wea,
        addra     => VMSME_L4PHIDn2_writeaddr,
        dina      => VMSME_L4PHIDn2_din,
        wea_out       => VMSME_L4PHIDn2_wea_delay,
        addra_out     => VMSME_L4PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L4PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L4PHIDn2_start
      );

    VMSME_L5PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L5PHIAn2_V_datatmp,
        dataout0 => VMSME_L5PHIAn2_AV_dout(0),
        dataout1 => VMSME_L5PHIAn2_AV_dout(1),
        dataout2 => VMSME_L5PHIAn2_AV_dout(2),
        dataout3 => VMSME_L5PHIAn2_AV_dout(3)
      );

    VMSME_L5PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L5PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L5PHIAn2_wea_delay,
        addra     => VMSME_L5PHIAn2_writeaddr_delay,
        dina      => VMSME_L5PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L5PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L5PHIAn2_AV_readaddr(3),VMSME_L5PHIAn2_AV_readaddr(2),VMSME_L5PHIAn2_AV_readaddr(1),VMSME_L5PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L5PHIAn2_V_datatmp,
        enb_nent  => VMSME_L5PHIAn2_enb_nent,
        addr_nent  => VMSME_L5PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L5PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L5PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L5PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L5PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L5PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L5PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L5PHIAn2_V_binmaskb
      );

    VMSME_L5PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L5PHIAn2_wea,
        addra     => VMSME_L5PHIAn2_writeaddr,
        dina      => VMSME_L5PHIAn2_din,
        wea_out       => VMSME_L5PHIAn2_wea_delay,
        addra_out     => VMSME_L5PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L5PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L5PHIAn2_start
      );

    VMSME_L5PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L5PHIBn2_V_datatmp,
        dataout0 => VMSME_L5PHIBn2_AV_dout(0),
        dataout1 => VMSME_L5PHIBn2_AV_dout(1),
        dataout2 => VMSME_L5PHIBn2_AV_dout(2),
        dataout3 => VMSME_L5PHIBn2_AV_dout(3)
      );

    VMSME_L5PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L5PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L5PHIBn2_wea_delay,
        addra     => VMSME_L5PHIBn2_writeaddr_delay,
        dina      => VMSME_L5PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L5PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L5PHIBn2_AV_readaddr(3),VMSME_L5PHIBn2_AV_readaddr(2),VMSME_L5PHIBn2_AV_readaddr(1),VMSME_L5PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L5PHIBn2_V_datatmp,
        enb_nent  => VMSME_L5PHIBn2_enb_nent,
        addr_nent  => VMSME_L5PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L5PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L5PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L5PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L5PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L5PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L5PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L5PHIBn2_V_binmaskb
      );

    VMSME_L5PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L5PHIBn2_wea,
        addra     => VMSME_L5PHIBn2_writeaddr,
        dina      => VMSME_L5PHIBn2_din,
        wea_out       => VMSME_L5PHIBn2_wea_delay,
        addra_out     => VMSME_L5PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L5PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L5PHIBn2_start
      );

    VMSME_L5PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L5PHICn2_V_datatmp,
        dataout0 => VMSME_L5PHICn2_AV_dout(0),
        dataout1 => VMSME_L5PHICn2_AV_dout(1),
        dataout2 => VMSME_L5PHICn2_AV_dout(2),
        dataout3 => VMSME_L5PHICn2_AV_dout(3)
      );

    VMSME_L5PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L5PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L5PHICn2_wea_delay,
        addra     => VMSME_L5PHICn2_writeaddr_delay,
        dina      => VMSME_L5PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L5PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L5PHICn2_AV_readaddr(3),VMSME_L5PHICn2_AV_readaddr(2),VMSME_L5PHICn2_AV_readaddr(1),VMSME_L5PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L5PHICn2_V_datatmp,
        enb_nent  => VMSME_L5PHICn2_enb_nent,
        addr_nent  => VMSME_L5PHICn2_V_addr_nent,
        dout_nent  => VMSME_L5PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L5PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L5PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L5PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L5PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L5PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L5PHICn2_V_binmaskb
      );

    VMSME_L5PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L5PHICn2_wea,
        addra     => VMSME_L5PHICn2_writeaddr,
        dina      => VMSME_L5PHICn2_din,
        wea_out       => VMSME_L5PHICn2_wea_delay,
        addra_out     => VMSME_L5PHICn2_writeaddr_delay,
        dina_out      => VMSME_L5PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L5PHICn2_start
      );

    VMSME_L5PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L5PHIDn2_V_datatmp,
        dataout0 => VMSME_L5PHIDn2_AV_dout(0),
        dataout1 => VMSME_L5PHIDn2_AV_dout(1),
        dataout2 => VMSME_L5PHIDn2_AV_dout(2),
        dataout3 => VMSME_L5PHIDn2_AV_dout(3)
      );

    VMSME_L5PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L5PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L5PHIDn2_wea_delay,
        addra     => VMSME_L5PHIDn2_writeaddr_delay,
        dina      => VMSME_L5PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L5PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L5PHIDn2_AV_readaddr(3),VMSME_L5PHIDn2_AV_readaddr(2),VMSME_L5PHIDn2_AV_readaddr(1),VMSME_L5PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L5PHIDn2_V_datatmp,
        enb_nent  => VMSME_L5PHIDn2_enb_nent,
        addr_nent  => VMSME_L5PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L5PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L5PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L5PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L5PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L5PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L5PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L5PHIDn2_V_binmaskb
      );

    VMSME_L5PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L5PHIDn2_wea,
        addra     => VMSME_L5PHIDn2_writeaddr,
        dina      => VMSME_L5PHIDn2_din,
        wea_out       => VMSME_L5PHIDn2_wea_delay,
        addra_out     => VMSME_L5PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L5PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L5PHIDn2_start
      );

    VMSME_L6PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L6PHIAn2_V_datatmp,
        dataout0 => VMSME_L6PHIAn2_AV_dout(0),
        dataout1 => VMSME_L6PHIAn2_AV_dout(1),
        dataout2 => VMSME_L6PHIAn2_AV_dout(2),
        dataout3 => VMSME_L6PHIAn2_AV_dout(3)
      );

    VMSME_L6PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L6PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L6PHIAn2_wea_delay,
        addra     => VMSME_L6PHIAn2_writeaddr_delay,
        dina      => VMSME_L6PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L6PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L6PHIAn2_AV_readaddr(3),VMSME_L6PHIAn2_AV_readaddr(2),VMSME_L6PHIAn2_AV_readaddr(1),VMSME_L6PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_L6PHIAn2_V_datatmp,
        enb_nent  => VMSME_L6PHIAn2_enb_nent,
        addr_nent  => VMSME_L6PHIAn2_V_addr_nent,
        dout_nent  => VMSME_L6PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_L6PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_L6PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_L6PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_L6PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L6PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L6PHIAn2_V_binmaskb
      );

    VMSME_L6PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L6PHIAn2_wea,
        addra     => VMSME_L6PHIAn2_writeaddr,
        dina      => VMSME_L6PHIAn2_din,
        wea_out       => VMSME_L6PHIAn2_wea_delay,
        addra_out     => VMSME_L6PHIAn2_writeaddr_delay,
        dina_out      => VMSME_L6PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_L6PHIAn2_start
      );

    VMSME_L6PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L6PHIBn2_V_datatmp,
        dataout0 => VMSME_L6PHIBn2_AV_dout(0),
        dataout1 => VMSME_L6PHIBn2_AV_dout(1),
        dataout2 => VMSME_L6PHIBn2_AV_dout(2),
        dataout3 => VMSME_L6PHIBn2_AV_dout(3)
      );

    VMSME_L6PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L6PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L6PHIBn2_wea_delay,
        addra     => VMSME_L6PHIBn2_writeaddr_delay,
        dina      => VMSME_L6PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L6PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L6PHIBn2_AV_readaddr(3),VMSME_L6PHIBn2_AV_readaddr(2),VMSME_L6PHIBn2_AV_readaddr(1),VMSME_L6PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_L6PHIBn2_V_datatmp,
        enb_nent  => VMSME_L6PHIBn2_enb_nent,
        addr_nent  => VMSME_L6PHIBn2_V_addr_nent,
        dout_nent  => VMSME_L6PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_L6PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_L6PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_L6PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_L6PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L6PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L6PHIBn2_V_binmaskb
      );

    VMSME_L6PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L6PHIBn2_wea,
        addra     => VMSME_L6PHIBn2_writeaddr,
        dina      => VMSME_L6PHIBn2_din,
        wea_out       => VMSME_L6PHIBn2_wea_delay,
        addra_out     => VMSME_L6PHIBn2_writeaddr_delay,
        dina_out      => VMSME_L6PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_L6PHIBn2_start
      );

    VMSME_L6PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L6PHICn2_V_datatmp,
        dataout0 => VMSME_L6PHICn2_AV_dout(0),
        dataout1 => VMSME_L6PHICn2_AV_dout(1),
        dataout2 => VMSME_L6PHICn2_AV_dout(2),
        dataout3 => VMSME_L6PHICn2_AV_dout(3)
      );

    VMSME_L6PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L6PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L6PHICn2_wea_delay,
        addra     => VMSME_L6PHICn2_writeaddr_delay,
        dina      => VMSME_L6PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L6PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L6PHICn2_AV_readaddr(3),VMSME_L6PHICn2_AV_readaddr(2),VMSME_L6PHICn2_AV_readaddr(1),VMSME_L6PHICn2_AV_readaddr(0)),
        doutb     => VMSME_L6PHICn2_V_datatmp,
        enb_nent  => VMSME_L6PHICn2_enb_nent,
        addr_nent  => VMSME_L6PHICn2_V_addr_nent,
        dout_nent  => VMSME_L6PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_L6PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_L6PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_L6PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_L6PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L6PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L6PHICn2_V_binmaskb
      );

    VMSME_L6PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L6PHICn2_wea,
        addra     => VMSME_L6PHICn2_writeaddr,
        dina      => VMSME_L6PHICn2_din,
        wea_out       => VMSME_L6PHICn2_wea_delay,
        addra_out     => VMSME_L6PHICn2_writeaddr_delay,
        dina_out      => VMSME_L6PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_L6PHICn2_start
      );

    VMSME_L6PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_L6PHIDn2_V_datatmp,
        dataout0 => VMSME_L6PHIDn2_AV_dout(0),
        dataout1 => VMSME_L6PHIDn2_AV_dout(1),
        dataout2 => VMSME_L6PHIDn2_AV_dout(2),
        dataout3 => VMSME_L6PHIDn2_AV_dout(3)
      );

    VMSME_L6PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_L6PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_L6PHIDn2_wea_delay,
        addra     => VMSME_L6PHIDn2_writeaddr_delay,
        dina      => VMSME_L6PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_L6PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_L6PHIDn2_AV_readaddr(3),VMSME_L6PHIDn2_AV_readaddr(2),VMSME_L6PHIDn2_AV_readaddr(1),VMSME_L6PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_L6PHIDn2_V_datatmp,
        enb_nent  => VMSME_L6PHIDn2_enb_nent,
        addr_nent  => VMSME_L6PHIDn2_V_addr_nent,
        dout_nent  => VMSME_L6PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_L6PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_L6PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_L6PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_L6PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_L6PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_L6PHIDn2_V_binmaskb
      );

    VMSME_L6PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_L6PHIDn2_wea,
        addra     => VMSME_L6PHIDn2_writeaddr,
        dina      => VMSME_L6PHIDn2_din,
        wea_out       => VMSME_L6PHIDn2_wea_delay,
        addra_out     => VMSME_L6PHIDn2_writeaddr_delay,
        dina_out      => VMSME_L6PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_L6PHIDn2_start
      );

    VMSME_D1PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D1PHIAn2_V_datatmp,
        dataout0 => VMSME_D1PHIAn2_AV_dout(0),
        dataout1 => VMSME_D1PHIAn2_AV_dout(1),
        dataout2 => VMSME_D1PHIAn2_AV_dout(2),
        dataout3 => VMSME_D1PHIAn2_AV_dout(3)
      );

    VMSME_D1PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D1PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D1PHIAn2_wea_delay,
        addra     => VMSME_D1PHIAn2_writeaddr_delay,
        dina      => VMSME_D1PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D1PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D1PHIAn2_AV_readaddr(3),VMSME_D1PHIAn2_AV_readaddr(2),VMSME_D1PHIAn2_AV_readaddr(1),VMSME_D1PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_D1PHIAn2_V_datatmp,
        enb_nent  => VMSME_D1PHIAn2_enb_nent,
        addr_nent  => VMSME_D1PHIAn2_V_addr_nent,
        dout_nent  => VMSME_D1PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_D1PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_D1PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_D1PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_D1PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D1PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D1PHIAn2_V_binmaskb
      );

    VMSME_D1PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D1PHIAn2_wea,
        addra     => VMSME_D1PHIAn2_writeaddr,
        dina      => VMSME_D1PHIAn2_din,
        wea_out       => VMSME_D1PHIAn2_wea_delay,
        addra_out     => VMSME_D1PHIAn2_writeaddr_delay,
        dina_out      => VMSME_D1PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_D1PHIAn2_start
      );

    VMSME_D1PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D1PHIBn2_V_datatmp,
        dataout0 => VMSME_D1PHIBn2_AV_dout(0),
        dataout1 => VMSME_D1PHIBn2_AV_dout(1),
        dataout2 => VMSME_D1PHIBn2_AV_dout(2),
        dataout3 => VMSME_D1PHIBn2_AV_dout(3)
      );

    VMSME_D1PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D1PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D1PHIBn2_wea_delay,
        addra     => VMSME_D1PHIBn2_writeaddr_delay,
        dina      => VMSME_D1PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D1PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D1PHIBn2_AV_readaddr(3),VMSME_D1PHIBn2_AV_readaddr(2),VMSME_D1PHIBn2_AV_readaddr(1),VMSME_D1PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_D1PHIBn2_V_datatmp,
        enb_nent  => VMSME_D1PHIBn2_enb_nent,
        addr_nent  => VMSME_D1PHIBn2_V_addr_nent,
        dout_nent  => VMSME_D1PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_D1PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_D1PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_D1PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_D1PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D1PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D1PHIBn2_V_binmaskb
      );

    VMSME_D1PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D1PHIBn2_wea,
        addra     => VMSME_D1PHIBn2_writeaddr,
        dina      => VMSME_D1PHIBn2_din,
        wea_out       => VMSME_D1PHIBn2_wea_delay,
        addra_out     => VMSME_D1PHIBn2_writeaddr_delay,
        dina_out      => VMSME_D1PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_D1PHIBn2_start
      );

    VMSME_D1PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D1PHICn2_V_datatmp,
        dataout0 => VMSME_D1PHICn2_AV_dout(0),
        dataout1 => VMSME_D1PHICn2_AV_dout(1),
        dataout2 => VMSME_D1PHICn2_AV_dout(2),
        dataout3 => VMSME_D1PHICn2_AV_dout(3)
      );

    VMSME_D1PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D1PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D1PHICn2_wea_delay,
        addra     => VMSME_D1PHICn2_writeaddr_delay,
        dina      => VMSME_D1PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D1PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D1PHICn2_AV_readaddr(3),VMSME_D1PHICn2_AV_readaddr(2),VMSME_D1PHICn2_AV_readaddr(1),VMSME_D1PHICn2_AV_readaddr(0)),
        doutb     => VMSME_D1PHICn2_V_datatmp,
        enb_nent  => VMSME_D1PHICn2_enb_nent,
        addr_nent  => VMSME_D1PHICn2_V_addr_nent,
        dout_nent  => VMSME_D1PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_D1PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_D1PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_D1PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_D1PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D1PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D1PHICn2_V_binmaskb
      );

    VMSME_D1PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D1PHICn2_wea,
        addra     => VMSME_D1PHICn2_writeaddr,
        dina      => VMSME_D1PHICn2_din,
        wea_out       => VMSME_D1PHICn2_wea_delay,
        addra_out     => VMSME_D1PHICn2_writeaddr_delay,
        dina_out      => VMSME_D1PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_D1PHICn2_start
      );

    VMSME_D1PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D1PHIDn2_V_datatmp,
        dataout0 => VMSME_D1PHIDn2_AV_dout(0),
        dataout1 => VMSME_D1PHIDn2_AV_dout(1),
        dataout2 => VMSME_D1PHIDn2_AV_dout(2),
        dataout3 => VMSME_D1PHIDn2_AV_dout(3)
      );

    VMSME_D1PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D1PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D1PHIDn2_wea_delay,
        addra     => VMSME_D1PHIDn2_writeaddr_delay,
        dina      => VMSME_D1PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D1PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D1PHIDn2_AV_readaddr(3),VMSME_D1PHIDn2_AV_readaddr(2),VMSME_D1PHIDn2_AV_readaddr(1),VMSME_D1PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_D1PHIDn2_V_datatmp,
        enb_nent  => VMSME_D1PHIDn2_enb_nent,
        addr_nent  => VMSME_D1PHIDn2_V_addr_nent,
        dout_nent  => VMSME_D1PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_D1PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_D1PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_D1PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_D1PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D1PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D1PHIDn2_V_binmaskb
      );

    VMSME_D1PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D1PHIDn2_wea,
        addra     => VMSME_D1PHIDn2_writeaddr,
        dina      => VMSME_D1PHIDn2_din,
        wea_out       => VMSME_D1PHIDn2_wea_delay,
        addra_out     => VMSME_D1PHIDn2_writeaddr_delay,
        dina_out      => VMSME_D1PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_D1PHIDn2_start
      );

    VMSME_D2PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D2PHIAn2_V_datatmp,
        dataout0 => VMSME_D2PHIAn2_AV_dout(0),
        dataout1 => VMSME_D2PHIAn2_AV_dout(1),
        dataout2 => VMSME_D2PHIAn2_AV_dout(2),
        dataout3 => VMSME_D2PHIAn2_AV_dout(3)
      );

    VMSME_D2PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D2PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D2PHIAn2_wea_delay,
        addra     => VMSME_D2PHIAn2_writeaddr_delay,
        dina      => VMSME_D2PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D2PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D2PHIAn2_AV_readaddr(3),VMSME_D2PHIAn2_AV_readaddr(2),VMSME_D2PHIAn2_AV_readaddr(1),VMSME_D2PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_D2PHIAn2_V_datatmp,
        enb_nent  => VMSME_D2PHIAn2_enb_nent,
        addr_nent  => VMSME_D2PHIAn2_V_addr_nent,
        dout_nent  => VMSME_D2PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_D2PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_D2PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_D2PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_D2PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D2PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D2PHIAn2_V_binmaskb
      );

    VMSME_D2PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D2PHIAn2_wea,
        addra     => VMSME_D2PHIAn2_writeaddr,
        dina      => VMSME_D2PHIAn2_din,
        wea_out       => VMSME_D2PHIAn2_wea_delay,
        addra_out     => VMSME_D2PHIAn2_writeaddr_delay,
        dina_out      => VMSME_D2PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_D2PHIAn2_start
      );

    VMSME_D2PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D2PHIBn2_V_datatmp,
        dataout0 => VMSME_D2PHIBn2_AV_dout(0),
        dataout1 => VMSME_D2PHIBn2_AV_dout(1),
        dataout2 => VMSME_D2PHIBn2_AV_dout(2),
        dataout3 => VMSME_D2PHIBn2_AV_dout(3)
      );

    VMSME_D2PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D2PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D2PHIBn2_wea_delay,
        addra     => VMSME_D2PHIBn2_writeaddr_delay,
        dina      => VMSME_D2PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D2PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D2PHIBn2_AV_readaddr(3),VMSME_D2PHIBn2_AV_readaddr(2),VMSME_D2PHIBn2_AV_readaddr(1),VMSME_D2PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_D2PHIBn2_V_datatmp,
        enb_nent  => VMSME_D2PHIBn2_enb_nent,
        addr_nent  => VMSME_D2PHIBn2_V_addr_nent,
        dout_nent  => VMSME_D2PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_D2PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_D2PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_D2PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_D2PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D2PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D2PHIBn2_V_binmaskb
      );

    VMSME_D2PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D2PHIBn2_wea,
        addra     => VMSME_D2PHIBn2_writeaddr,
        dina      => VMSME_D2PHIBn2_din,
        wea_out       => VMSME_D2PHIBn2_wea_delay,
        addra_out     => VMSME_D2PHIBn2_writeaddr_delay,
        dina_out      => VMSME_D2PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_D2PHIBn2_start
      );

    VMSME_D2PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D2PHICn2_V_datatmp,
        dataout0 => VMSME_D2PHICn2_AV_dout(0),
        dataout1 => VMSME_D2PHICn2_AV_dout(1),
        dataout2 => VMSME_D2PHICn2_AV_dout(2),
        dataout3 => VMSME_D2PHICn2_AV_dout(3)
      );

    VMSME_D2PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D2PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D2PHICn2_wea_delay,
        addra     => VMSME_D2PHICn2_writeaddr_delay,
        dina      => VMSME_D2PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D2PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D2PHICn2_AV_readaddr(3),VMSME_D2PHICn2_AV_readaddr(2),VMSME_D2PHICn2_AV_readaddr(1),VMSME_D2PHICn2_AV_readaddr(0)),
        doutb     => VMSME_D2PHICn2_V_datatmp,
        enb_nent  => VMSME_D2PHICn2_enb_nent,
        addr_nent  => VMSME_D2PHICn2_V_addr_nent,
        dout_nent  => VMSME_D2PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_D2PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_D2PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_D2PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_D2PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D2PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D2PHICn2_V_binmaskb
      );

    VMSME_D2PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D2PHICn2_wea,
        addra     => VMSME_D2PHICn2_writeaddr,
        dina      => VMSME_D2PHICn2_din,
        wea_out       => VMSME_D2PHICn2_wea_delay,
        addra_out     => VMSME_D2PHICn2_writeaddr_delay,
        dina_out      => VMSME_D2PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_D2PHICn2_start
      );

    VMSME_D2PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D2PHIDn2_V_datatmp,
        dataout0 => VMSME_D2PHIDn2_AV_dout(0),
        dataout1 => VMSME_D2PHIDn2_AV_dout(1),
        dataout2 => VMSME_D2PHIDn2_AV_dout(2),
        dataout3 => VMSME_D2PHIDn2_AV_dout(3)
      );

    VMSME_D2PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D2PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D2PHIDn2_wea_delay,
        addra     => VMSME_D2PHIDn2_writeaddr_delay,
        dina      => VMSME_D2PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D2PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D2PHIDn2_AV_readaddr(3),VMSME_D2PHIDn2_AV_readaddr(2),VMSME_D2PHIDn2_AV_readaddr(1),VMSME_D2PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_D2PHIDn2_V_datatmp,
        enb_nent  => VMSME_D2PHIDn2_enb_nent,
        addr_nent  => VMSME_D2PHIDn2_V_addr_nent,
        dout_nent  => VMSME_D2PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_D2PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_D2PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_D2PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_D2PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D2PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D2PHIDn2_V_binmaskb
      );

    VMSME_D2PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D2PHIDn2_wea,
        addra     => VMSME_D2PHIDn2_writeaddr,
        dina      => VMSME_D2PHIDn2_din,
        wea_out       => VMSME_D2PHIDn2_wea_delay,
        addra_out     => VMSME_D2PHIDn2_writeaddr_delay,
        dina_out      => VMSME_D2PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_D2PHIDn2_start
      );

    VMSME_D3PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D3PHIAn2_V_datatmp,
        dataout0 => VMSME_D3PHIAn2_AV_dout(0),
        dataout1 => VMSME_D3PHIAn2_AV_dout(1),
        dataout2 => VMSME_D3PHIAn2_AV_dout(2),
        dataout3 => VMSME_D3PHIAn2_AV_dout(3)
      );

    VMSME_D3PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D3PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D3PHIAn2_wea_delay,
        addra     => VMSME_D3PHIAn2_writeaddr_delay,
        dina      => VMSME_D3PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D3PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D3PHIAn2_AV_readaddr(3),VMSME_D3PHIAn2_AV_readaddr(2),VMSME_D3PHIAn2_AV_readaddr(1),VMSME_D3PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_D3PHIAn2_V_datatmp,
        enb_nent  => VMSME_D3PHIAn2_enb_nent,
        addr_nent  => VMSME_D3PHIAn2_V_addr_nent,
        dout_nent  => VMSME_D3PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_D3PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_D3PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_D3PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_D3PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D3PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D3PHIAn2_V_binmaskb
      );

    VMSME_D3PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D3PHIAn2_wea,
        addra     => VMSME_D3PHIAn2_writeaddr,
        dina      => VMSME_D3PHIAn2_din,
        wea_out       => VMSME_D3PHIAn2_wea_delay,
        addra_out     => VMSME_D3PHIAn2_writeaddr_delay,
        dina_out      => VMSME_D3PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_D3PHIAn2_start
      );

    VMSME_D3PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D3PHIBn2_V_datatmp,
        dataout0 => VMSME_D3PHIBn2_AV_dout(0),
        dataout1 => VMSME_D3PHIBn2_AV_dout(1),
        dataout2 => VMSME_D3PHIBn2_AV_dout(2),
        dataout3 => VMSME_D3PHIBn2_AV_dout(3)
      );

    VMSME_D3PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D3PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D3PHIBn2_wea_delay,
        addra     => VMSME_D3PHIBn2_writeaddr_delay,
        dina      => VMSME_D3PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D3PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D3PHIBn2_AV_readaddr(3),VMSME_D3PHIBn2_AV_readaddr(2),VMSME_D3PHIBn2_AV_readaddr(1),VMSME_D3PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_D3PHIBn2_V_datatmp,
        enb_nent  => VMSME_D3PHIBn2_enb_nent,
        addr_nent  => VMSME_D3PHIBn2_V_addr_nent,
        dout_nent  => VMSME_D3PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_D3PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_D3PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_D3PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_D3PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D3PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D3PHIBn2_V_binmaskb
      );

    VMSME_D3PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D3PHIBn2_wea,
        addra     => VMSME_D3PHIBn2_writeaddr,
        dina      => VMSME_D3PHIBn2_din,
        wea_out       => VMSME_D3PHIBn2_wea_delay,
        addra_out     => VMSME_D3PHIBn2_writeaddr_delay,
        dina_out      => VMSME_D3PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_D3PHIBn2_start
      );

    VMSME_D3PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D3PHICn2_V_datatmp,
        dataout0 => VMSME_D3PHICn2_AV_dout(0),
        dataout1 => VMSME_D3PHICn2_AV_dout(1),
        dataout2 => VMSME_D3PHICn2_AV_dout(2),
        dataout3 => VMSME_D3PHICn2_AV_dout(3)
      );

    VMSME_D3PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D3PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D3PHICn2_wea_delay,
        addra     => VMSME_D3PHICn2_writeaddr_delay,
        dina      => VMSME_D3PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D3PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D3PHICn2_AV_readaddr(3),VMSME_D3PHICn2_AV_readaddr(2),VMSME_D3PHICn2_AV_readaddr(1),VMSME_D3PHICn2_AV_readaddr(0)),
        doutb     => VMSME_D3PHICn2_V_datatmp,
        enb_nent  => VMSME_D3PHICn2_enb_nent,
        addr_nent  => VMSME_D3PHICn2_V_addr_nent,
        dout_nent  => VMSME_D3PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_D3PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_D3PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_D3PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_D3PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D3PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D3PHICn2_V_binmaskb
      );

    VMSME_D3PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D3PHICn2_wea,
        addra     => VMSME_D3PHICn2_writeaddr,
        dina      => VMSME_D3PHICn2_din,
        wea_out       => VMSME_D3PHICn2_wea_delay,
        addra_out     => VMSME_D3PHICn2_writeaddr_delay,
        dina_out      => VMSME_D3PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_D3PHICn2_start
      );

    VMSME_D3PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D3PHIDn2_V_datatmp,
        dataout0 => VMSME_D3PHIDn2_AV_dout(0),
        dataout1 => VMSME_D3PHIDn2_AV_dout(1),
        dataout2 => VMSME_D3PHIDn2_AV_dout(2),
        dataout3 => VMSME_D3PHIDn2_AV_dout(3)
      );

    VMSME_D3PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D3PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D3PHIDn2_wea_delay,
        addra     => VMSME_D3PHIDn2_writeaddr_delay,
        dina      => VMSME_D3PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D3PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D3PHIDn2_AV_readaddr(3),VMSME_D3PHIDn2_AV_readaddr(2),VMSME_D3PHIDn2_AV_readaddr(1),VMSME_D3PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_D3PHIDn2_V_datatmp,
        enb_nent  => VMSME_D3PHIDn2_enb_nent,
        addr_nent  => VMSME_D3PHIDn2_V_addr_nent,
        dout_nent  => VMSME_D3PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_D3PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_D3PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_D3PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_D3PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D3PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D3PHIDn2_V_binmaskb
      );

    VMSME_D3PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D3PHIDn2_wea,
        addra     => VMSME_D3PHIDn2_writeaddr,
        dina      => VMSME_D3PHIDn2_din,
        wea_out       => VMSME_D3PHIDn2_wea_delay,
        addra_out     => VMSME_D3PHIDn2_writeaddr_delay,
        dina_out      => VMSME_D3PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_D3PHIDn2_start
      );

    VMSME_D4PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D4PHIAn2_V_datatmp,
        dataout0 => VMSME_D4PHIAn2_AV_dout(0),
        dataout1 => VMSME_D4PHIAn2_AV_dout(1),
        dataout2 => VMSME_D4PHIAn2_AV_dout(2),
        dataout3 => VMSME_D4PHIAn2_AV_dout(3)
      );

    VMSME_D4PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D4PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D4PHIAn2_wea_delay,
        addra     => VMSME_D4PHIAn2_writeaddr_delay,
        dina      => VMSME_D4PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D4PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D4PHIAn2_AV_readaddr(3),VMSME_D4PHIAn2_AV_readaddr(2),VMSME_D4PHIAn2_AV_readaddr(1),VMSME_D4PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_D4PHIAn2_V_datatmp,
        enb_nent  => VMSME_D4PHIAn2_enb_nent,
        addr_nent  => VMSME_D4PHIAn2_V_addr_nent,
        dout_nent  => VMSME_D4PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_D4PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_D4PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_D4PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_D4PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D4PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D4PHIAn2_V_binmaskb
      );

    VMSME_D4PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D4PHIAn2_wea,
        addra     => VMSME_D4PHIAn2_writeaddr,
        dina      => VMSME_D4PHIAn2_din,
        wea_out       => VMSME_D4PHIAn2_wea_delay,
        addra_out     => VMSME_D4PHIAn2_writeaddr_delay,
        dina_out      => VMSME_D4PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_D4PHIAn2_start
      );

    VMSME_D4PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D4PHIBn2_V_datatmp,
        dataout0 => VMSME_D4PHIBn2_AV_dout(0),
        dataout1 => VMSME_D4PHIBn2_AV_dout(1),
        dataout2 => VMSME_D4PHIBn2_AV_dout(2),
        dataout3 => VMSME_D4PHIBn2_AV_dout(3)
      );

    VMSME_D4PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D4PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D4PHIBn2_wea_delay,
        addra     => VMSME_D4PHIBn2_writeaddr_delay,
        dina      => VMSME_D4PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D4PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D4PHIBn2_AV_readaddr(3),VMSME_D4PHIBn2_AV_readaddr(2),VMSME_D4PHIBn2_AV_readaddr(1),VMSME_D4PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_D4PHIBn2_V_datatmp,
        enb_nent  => VMSME_D4PHIBn2_enb_nent,
        addr_nent  => VMSME_D4PHIBn2_V_addr_nent,
        dout_nent  => VMSME_D4PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_D4PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_D4PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_D4PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_D4PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D4PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D4PHIBn2_V_binmaskb
      );

    VMSME_D4PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D4PHIBn2_wea,
        addra     => VMSME_D4PHIBn2_writeaddr,
        dina      => VMSME_D4PHIBn2_din,
        wea_out       => VMSME_D4PHIBn2_wea_delay,
        addra_out     => VMSME_D4PHIBn2_writeaddr_delay,
        dina_out      => VMSME_D4PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_D4PHIBn2_start
      );

    VMSME_D4PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D4PHICn2_V_datatmp,
        dataout0 => VMSME_D4PHICn2_AV_dout(0),
        dataout1 => VMSME_D4PHICn2_AV_dout(1),
        dataout2 => VMSME_D4PHICn2_AV_dout(2),
        dataout3 => VMSME_D4PHICn2_AV_dout(3)
      );

    VMSME_D4PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D4PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D4PHICn2_wea_delay,
        addra     => VMSME_D4PHICn2_writeaddr_delay,
        dina      => VMSME_D4PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D4PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D4PHICn2_AV_readaddr(3),VMSME_D4PHICn2_AV_readaddr(2),VMSME_D4PHICn2_AV_readaddr(1),VMSME_D4PHICn2_AV_readaddr(0)),
        doutb     => VMSME_D4PHICn2_V_datatmp,
        enb_nent  => VMSME_D4PHICn2_enb_nent,
        addr_nent  => VMSME_D4PHICn2_V_addr_nent,
        dout_nent  => VMSME_D4PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_D4PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_D4PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_D4PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_D4PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D4PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D4PHICn2_V_binmaskb
      );

    VMSME_D4PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D4PHICn2_wea,
        addra     => VMSME_D4PHICn2_writeaddr,
        dina      => VMSME_D4PHICn2_din,
        wea_out       => VMSME_D4PHICn2_wea_delay,
        addra_out     => VMSME_D4PHICn2_writeaddr_delay,
        dina_out      => VMSME_D4PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_D4PHICn2_start
      );

    VMSME_D4PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D4PHIDn2_V_datatmp,
        dataout0 => VMSME_D4PHIDn2_AV_dout(0),
        dataout1 => VMSME_D4PHIDn2_AV_dout(1),
        dataout2 => VMSME_D4PHIDn2_AV_dout(2),
        dataout3 => VMSME_D4PHIDn2_AV_dout(3)
      );

    VMSME_D4PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D4PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D4PHIDn2_wea_delay,
        addra     => VMSME_D4PHIDn2_writeaddr_delay,
        dina      => VMSME_D4PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D4PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D4PHIDn2_AV_readaddr(3),VMSME_D4PHIDn2_AV_readaddr(2),VMSME_D4PHIDn2_AV_readaddr(1),VMSME_D4PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_D4PHIDn2_V_datatmp,
        enb_nent  => VMSME_D4PHIDn2_enb_nent,
        addr_nent  => VMSME_D4PHIDn2_V_addr_nent,
        dout_nent  => VMSME_D4PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_D4PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_D4PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_D4PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_D4PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D4PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D4PHIDn2_V_binmaskb
      );

    VMSME_D4PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D4PHIDn2_wea,
        addra     => VMSME_D4PHIDn2_writeaddr,
        dina      => VMSME_D4PHIDn2_din,
        wea_out       => VMSME_D4PHIDn2_wea_delay,
        addra_out     => VMSME_D4PHIDn2_writeaddr_delay,
        dina_out      => VMSME_D4PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_D4PHIDn2_start
      );

    VMSME_D5PHIAn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D5PHIAn2_V_datatmp,
        dataout0 => VMSME_D5PHIAn2_AV_dout(0),
        dataout1 => VMSME_D5PHIAn2_AV_dout(1),
        dataout2 => VMSME_D5PHIAn2_AV_dout(2),
        dataout3 => VMSME_D5PHIAn2_AV_dout(3)
      );

    VMSME_D5PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D5PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D5PHIAn2_wea_delay,
        addra     => VMSME_D5PHIAn2_writeaddr_delay,
        dina      => VMSME_D5PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D5PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D5PHIAn2_AV_readaddr(3),VMSME_D5PHIAn2_AV_readaddr(2),VMSME_D5PHIAn2_AV_readaddr(1),VMSME_D5PHIAn2_AV_readaddr(0)),
        doutb     => VMSME_D5PHIAn2_V_datatmp,
        enb_nent  => VMSME_D5PHIAn2_enb_nent,
        addr_nent  => VMSME_D5PHIAn2_V_addr_nent,
        dout_nent  => VMSME_D5PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSME_D5PHIAn2_enb_binmaska,
        addr_binmaska  => VMSME_D5PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSME_D5PHIAn2_V_binmaska,
        enb_binmaskb  => VMSME_D5PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D5PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D5PHIAn2_V_binmaskb
      );

    VMSME_D5PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D5PHIAn2_wea,
        addra     => VMSME_D5PHIAn2_writeaddr,
        dina      => VMSME_D5PHIAn2_din,
        wea_out       => VMSME_D5PHIAn2_wea_delay,
        addra_out     => VMSME_D5PHIAn2_writeaddr_delay,
        dina_out      => VMSME_D5PHIAn2_din_delay,
        done       => PC_done,
        start      => VMSME_D5PHIAn2_start
      );

    VMSME_D5PHIBn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D5PHIBn2_V_datatmp,
        dataout0 => VMSME_D5PHIBn2_AV_dout(0),
        dataout1 => VMSME_D5PHIBn2_AV_dout(1),
        dataout2 => VMSME_D5PHIBn2_AV_dout(2),
        dataout3 => VMSME_D5PHIBn2_AV_dout(3)
      );

    VMSME_D5PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D5PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D5PHIBn2_wea_delay,
        addra     => VMSME_D5PHIBn2_writeaddr_delay,
        dina      => VMSME_D5PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D5PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D5PHIBn2_AV_readaddr(3),VMSME_D5PHIBn2_AV_readaddr(2),VMSME_D5PHIBn2_AV_readaddr(1),VMSME_D5PHIBn2_AV_readaddr(0)),
        doutb     => VMSME_D5PHIBn2_V_datatmp,
        enb_nent  => VMSME_D5PHIBn2_enb_nent,
        addr_nent  => VMSME_D5PHIBn2_V_addr_nent,
        dout_nent  => VMSME_D5PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSME_D5PHIBn2_enb_binmaska,
        addr_binmaska  => VMSME_D5PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSME_D5PHIBn2_V_binmaska,
        enb_binmaskb  => VMSME_D5PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D5PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D5PHIBn2_V_binmaskb
      );

    VMSME_D5PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D5PHIBn2_wea,
        addra     => VMSME_D5PHIBn2_writeaddr,
        dina      => VMSME_D5PHIBn2_din,
        wea_out       => VMSME_D5PHIBn2_wea_delay,
        addra_out     => VMSME_D5PHIBn2_writeaddr_delay,
        dina_out      => VMSME_D5PHIBn2_din_delay,
        done       => PC_done,
        start      => VMSME_D5PHIBn2_start
      );

    VMSME_D5PHICn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D5PHICn2_V_datatmp,
        dataout0 => VMSME_D5PHICn2_AV_dout(0),
        dataout1 => VMSME_D5PHICn2_AV_dout(1),
        dataout2 => VMSME_D5PHICn2_AV_dout(2),
        dataout3 => VMSME_D5PHICn2_AV_dout(3)
      );

    VMSME_D5PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D5PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D5PHICn2_wea_delay,
        addra     => VMSME_D5PHICn2_writeaddr_delay,
        dina      => VMSME_D5PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D5PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D5PHICn2_AV_readaddr(3),VMSME_D5PHICn2_AV_readaddr(2),VMSME_D5PHICn2_AV_readaddr(1),VMSME_D5PHICn2_AV_readaddr(0)),
        doutb     => VMSME_D5PHICn2_V_datatmp,
        enb_nent  => VMSME_D5PHICn2_enb_nent,
        addr_nent  => VMSME_D5PHICn2_V_addr_nent,
        dout_nent  => VMSME_D5PHICn2_AV_dout_nent,
        enb_binmaska  => VMSME_D5PHICn2_enb_binmaska,
        addr_binmaska  => VMSME_D5PHICn2_V_addr_binmaska,
        binmaska_o  => VMSME_D5PHICn2_V_binmaska,
        enb_binmaskb  => VMSME_D5PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D5PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D5PHICn2_V_binmaskb
      );

    VMSME_D5PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D5PHICn2_wea,
        addra     => VMSME_D5PHICn2_writeaddr,
        dina      => VMSME_D5PHICn2_din,
        wea_out       => VMSME_D5PHICn2_wea_delay,
        addra_out     => VMSME_D5PHICn2_writeaddr_delay,
        dina_out      => VMSME_D5PHICn2_din_delay,
        done       => PC_done,
        start      => VMSME_D5PHICn2_start
      );

    VMSME_D5PHIDn2_dataformat : entity work.vmstub17dout4
      port map (
        datain => VMSME_D5PHIDn2_V_datatmp,
        dataout0 => VMSME_D5PHIDn2_AV_dout(0),
        dataout1 => VMSME_D5PHIDn2_AV_dout(1),
        dataout2 => VMSME_D5PHIDn2_AV_dout(2),
        dataout3 => VMSME_D5PHIDn2_AV_dout(3)
      );

    VMSME_D5PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSME_D5PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 16,
        NUM_COPY        => 4
      )
      port map (
        clka      => clk,
        wea       => VMSME_D5PHIDn2_wea_delay,
        addra     => VMSME_D5PHIDn2_writeaddr_delay,
        dina      => VMSME_D5PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSME_D5PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSME_D5PHIDn2_AV_readaddr(3),VMSME_D5PHIDn2_AV_readaddr(2),VMSME_D5PHIDn2_AV_readaddr(1),VMSME_D5PHIDn2_AV_readaddr(0)),
        doutb     => VMSME_D5PHIDn2_V_datatmp,
        enb_nent  => VMSME_D5PHIDn2_enb_nent,
        addr_nent  => VMSME_D5PHIDn2_V_addr_nent,
        dout_nent  => VMSME_D5PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSME_D5PHIDn2_enb_binmaska,
        addr_binmaska  => VMSME_D5PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSME_D5PHIDn2_V_binmaska,
        enb_binmaskb  => VMSME_D5PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSME_D5PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSME_D5PHIDn2_V_binmaskb
      );

    VMSME_D5PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSME_D5PHIDn2_wea,
        addra     => VMSME_D5PHIDn2_writeaddr,
        dina      => VMSME_D5PHIDn2_din,
        wea_out       => VMSME_D5PHIDn2_wea_delay,
        addra_out     => VMSME_D5PHIDn2_writeaddr_delay,
        dina_out      => VMSME_D5PHIDn2_din_delay,
        done       => PC_done,
        start      => VMSME_D5PHIDn2_start
      );

    MPAR_L1L2ABCin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2ABCin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2ABCin_wea_delay,
        addra     => MPAR_L1L2ABCin_writeaddr_delay,
        dina      => MPAR_L1L2ABCin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2ABCin_V_readaddr,
        doutb     => MPAR_L1L2ABCin_V_dout,
        sync_nent => MPAR_L1L2ABCin_start,
        nent_o    => MPAR_L1L2ABCin_AV_dout_nent,
        mask_o    => MPAR_L1L2ABCin_AV_dout_mask
      );

    MPAR_L1L2ABCin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2ABCin_wea,
        addra     => MPAR_L1L2ABCin_writeaddr,
        dina      => MPAR_L1L2ABCin_din,
        wea_out       => MPAR_L1L2ABCin_wea_delay,
        addra_out     => MPAR_L1L2ABCin_writeaddr_delay,
        dina_out      => MPAR_L1L2ABCin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2ABCin_start
      );

    MPAR_L1L2DEin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2DEin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2DEin_wea_delay,
        addra     => MPAR_L1L2DEin_writeaddr_delay,
        dina      => MPAR_L1L2DEin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2DEin_V_readaddr,
        doutb     => MPAR_L1L2DEin_V_dout,
        sync_nent => MPAR_L1L2DEin_start,
        nent_o    => MPAR_L1L2DEin_AV_dout_nent,
        mask_o    => MPAR_L1L2DEin_AV_dout_mask
      );

    MPAR_L1L2DEin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2DEin_wea,
        addra     => MPAR_L1L2DEin_writeaddr,
        dina      => MPAR_L1L2DEin_din,
        wea_out       => MPAR_L1L2DEin_wea_delay,
        addra_out     => MPAR_L1L2DEin_writeaddr_delay,
        dina_out      => MPAR_L1L2DEin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2DEin_start
      );

    MPAR_L1L2Fin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2Fin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2Fin_wea_delay,
        addra     => MPAR_L1L2Fin_writeaddr_delay,
        dina      => MPAR_L1L2Fin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2Fin_V_readaddr,
        doutb     => MPAR_L1L2Fin_V_dout,
        sync_nent => MPAR_L1L2Fin_start,
        nent_o    => MPAR_L1L2Fin_AV_dout_nent,
        mask_o    => MPAR_L1L2Fin_AV_dout_mask
      );

    MPAR_L1L2Fin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2Fin_wea,
        addra     => MPAR_L1L2Fin_writeaddr,
        dina      => MPAR_L1L2Fin_din,
        wea_out       => MPAR_L1L2Fin_wea_delay,
        addra_out     => MPAR_L1L2Fin_writeaddr_delay,
        dina_out      => MPAR_L1L2Fin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2Fin_start
      );

    MPAR_L1L2Gin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2Gin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2Gin_wea_delay,
        addra     => MPAR_L1L2Gin_writeaddr_delay,
        dina      => MPAR_L1L2Gin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2Gin_V_readaddr,
        doutb     => MPAR_L1L2Gin_V_dout,
        sync_nent => MPAR_L1L2Gin_start,
        nent_o    => MPAR_L1L2Gin_AV_dout_nent,
        mask_o    => MPAR_L1L2Gin_AV_dout_mask
      );

    MPAR_L1L2Gin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2Gin_wea,
        addra     => MPAR_L1L2Gin_writeaddr,
        dina      => MPAR_L1L2Gin_din,
        wea_out       => MPAR_L1L2Gin_wea_delay,
        addra_out     => MPAR_L1L2Gin_writeaddr_delay,
        dina_out      => MPAR_L1L2Gin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2Gin_start
      );

    MPAR_L1L2HIin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2HIin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2HIin_wea_delay,
        addra     => MPAR_L1L2HIin_writeaddr_delay,
        dina      => MPAR_L1L2HIin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2HIin_V_readaddr,
        doutb     => MPAR_L1L2HIin_V_dout,
        sync_nent => MPAR_L1L2HIin_start,
        nent_o    => MPAR_L1L2HIin_AV_dout_nent,
        mask_o    => MPAR_L1L2HIin_AV_dout_mask
      );

    MPAR_L1L2HIin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2HIin_wea,
        addra     => MPAR_L1L2HIin_writeaddr,
        dina      => MPAR_L1L2HIin_din,
        wea_out       => MPAR_L1L2HIin_wea_delay,
        addra_out     => MPAR_L1L2HIin_writeaddr_delay,
        dina_out      => MPAR_L1L2HIin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2HIin_start
      );

    MPAR_L1L2JKLin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2JKLin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2JKLin_wea_delay,
        addra     => MPAR_L1L2JKLin_writeaddr_delay,
        dina      => MPAR_L1L2JKLin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2JKLin_V_readaddr,
        doutb     => MPAR_L1L2JKLin_V_dout,
        sync_nent => MPAR_L1L2JKLin_start,
        nent_o    => MPAR_L1L2JKLin_AV_dout_nent,
        mask_o    => MPAR_L1L2JKLin_AV_dout_mask
      );

    MPAR_L1L2JKLin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2JKLin_wea,
        addra     => MPAR_L1L2JKLin_writeaddr,
        dina      => MPAR_L1L2JKLin_din,
        wea_out       => MPAR_L1L2JKLin_wea_delay,
        addra_out     => MPAR_L1L2JKLin_writeaddr_delay,
        dina_out      => MPAR_L1L2JKLin_din_delay,
        done       => PC_start,
        start      => MPAR_L1L2JKLin_start
      );

    MPAR_L2L3ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L2L3ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L2L3ABCDin_wea_delay,
        addra     => MPAR_L2L3ABCDin_writeaddr_delay,
        dina      => MPAR_L2L3ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L2L3ABCDin_V_readaddr,
        doutb     => MPAR_L2L3ABCDin_V_dout,
        sync_nent => MPAR_L2L3ABCDin_start,
        nent_o    => MPAR_L2L3ABCDin_AV_dout_nent,
        mask_o    => MPAR_L2L3ABCDin_AV_dout_mask
      );

    MPAR_L2L3ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L2L3ABCDin_wea,
        addra     => MPAR_L2L3ABCDin_writeaddr,
        dina      => MPAR_L2L3ABCDin_din,
        wea_out       => MPAR_L2L3ABCDin_wea_delay,
        addra_out     => MPAR_L2L3ABCDin_writeaddr_delay,
        dina_out      => MPAR_L2L3ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_L2L3ABCDin_start
      );

    MPAR_L3L4ABin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L3L4ABin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L3L4ABin_wea_delay,
        addra     => MPAR_L3L4ABin_writeaddr_delay,
        dina      => MPAR_L3L4ABin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L3L4ABin_V_readaddr,
        doutb     => MPAR_L3L4ABin_V_dout,
        sync_nent => MPAR_L3L4ABin_start,
        nent_o    => MPAR_L3L4ABin_AV_dout_nent,
        mask_o    => MPAR_L3L4ABin_AV_dout_mask
      );

    MPAR_L3L4ABin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L3L4ABin_wea,
        addra     => MPAR_L3L4ABin_writeaddr,
        dina      => MPAR_L3L4ABin_din,
        wea_out       => MPAR_L3L4ABin_wea_delay,
        addra_out     => MPAR_L3L4ABin_writeaddr_delay,
        dina_out      => MPAR_L3L4ABin_din_delay,
        done       => PC_start,
        start      => MPAR_L3L4ABin_start
      );

    MPAR_L3L4CDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L3L4CDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L3L4CDin_wea_delay,
        addra     => MPAR_L3L4CDin_writeaddr_delay,
        dina      => MPAR_L3L4CDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L3L4CDin_V_readaddr,
        doutb     => MPAR_L3L4CDin_V_dout,
        sync_nent => MPAR_L3L4CDin_start,
        nent_o    => MPAR_L3L4CDin_AV_dout_nent,
        mask_o    => MPAR_L3L4CDin_AV_dout_mask
      );

    MPAR_L3L4CDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L3L4CDin_wea,
        addra     => MPAR_L3L4CDin_writeaddr,
        dina      => MPAR_L3L4CDin_din,
        wea_out       => MPAR_L3L4CDin_wea_delay,
        addra_out     => MPAR_L3L4CDin_writeaddr_delay,
        dina_out      => MPAR_L3L4CDin_din_delay,
        done       => PC_start,
        start      => MPAR_L3L4CDin_start
      );

    MPAR_L5L6ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L5L6ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L5L6ABCDin_wea_delay,
        addra     => MPAR_L5L6ABCDin_writeaddr_delay,
        dina      => MPAR_L5L6ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L5L6ABCDin_V_readaddr,
        doutb     => MPAR_L5L6ABCDin_V_dout,
        sync_nent => MPAR_L5L6ABCDin_start,
        nent_o    => MPAR_L5L6ABCDin_AV_dout_nent,
        mask_o    => MPAR_L5L6ABCDin_AV_dout_mask
      );

    MPAR_L5L6ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L5L6ABCDin_wea,
        addra     => MPAR_L5L6ABCDin_writeaddr,
        dina      => MPAR_L5L6ABCDin_din,
        wea_out       => MPAR_L5L6ABCDin_wea_delay,
        addra_out     => MPAR_L5L6ABCDin_writeaddr_delay,
        dina_out      => MPAR_L5L6ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_L5L6ABCDin_start
      );

    MPAR_D1D2ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_D1D2ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_D1D2ABCDin_wea_delay,
        addra     => MPAR_D1D2ABCDin_writeaddr_delay,
        dina      => MPAR_D1D2ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_D1D2ABCDin_V_readaddr,
        doutb     => MPAR_D1D2ABCDin_V_dout,
        sync_nent => MPAR_D1D2ABCDin_start,
        nent_o    => MPAR_D1D2ABCDin_AV_dout_nent,
        mask_o    => MPAR_D1D2ABCDin_AV_dout_mask
      );

    MPAR_D1D2ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_D1D2ABCDin_wea,
        addra     => MPAR_D1D2ABCDin_writeaddr,
        dina      => MPAR_D1D2ABCDin_din,
        wea_out       => MPAR_D1D2ABCDin_wea_delay,
        addra_out     => MPAR_D1D2ABCDin_writeaddr_delay,
        dina_out      => MPAR_D1D2ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_D1D2ABCDin_start
      );

    MPAR_D3D4ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_D3D4ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_D3D4ABCDin_wea_delay,
        addra     => MPAR_D3D4ABCDin_writeaddr_delay,
        dina      => MPAR_D3D4ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_D3D4ABCDin_V_readaddr,
        doutb     => MPAR_D3D4ABCDin_V_dout,
        sync_nent => MPAR_D3D4ABCDin_start,
        nent_o    => MPAR_D3D4ABCDin_AV_dout_nent,
        mask_o    => MPAR_D3D4ABCDin_AV_dout_mask
      );

    MPAR_D3D4ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_D3D4ABCDin_wea,
        addra     => MPAR_D3D4ABCDin_writeaddr,
        dina      => MPAR_D3D4ABCDin_din,
        wea_out       => MPAR_D3D4ABCDin_wea_delay,
        addra_out     => MPAR_D3D4ABCDin_writeaddr_delay,
        dina_out      => MPAR_D3D4ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_D3D4ABCDin_start
      );

    MPAR_L1D1ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1D1ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1D1ABCDin_wea_delay,
        addra     => MPAR_L1D1ABCDin_writeaddr_delay,
        dina      => MPAR_L1D1ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1D1ABCDin_V_readaddr,
        doutb     => MPAR_L1D1ABCDin_V_dout,
        sync_nent => MPAR_L1D1ABCDin_start,
        nent_o    => MPAR_L1D1ABCDin_AV_dout_nent,
        mask_o    => MPAR_L1D1ABCDin_AV_dout_mask
      );

    MPAR_L1D1ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1D1ABCDin_wea,
        addra     => MPAR_L1D1ABCDin_writeaddr,
        dina      => MPAR_L1D1ABCDin_din,
        wea_out       => MPAR_L1D1ABCDin_wea_delay,
        addra_out     => MPAR_L1D1ABCDin_writeaddr_delay,
        dina_out      => MPAR_L1D1ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_L1D1ABCDin_start
      );

    MPAR_L1D1EFGHin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1D1EFGHin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1D1EFGHin_wea_delay,
        addra     => MPAR_L1D1EFGHin_writeaddr_delay,
        dina      => MPAR_L1D1EFGHin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1D1EFGHin_V_readaddr,
        doutb     => MPAR_L1D1EFGHin_V_dout,
        sync_nent => MPAR_L1D1EFGHin_start,
        nent_o    => MPAR_L1D1EFGHin_AV_dout_nent,
        mask_o    => MPAR_L1D1EFGHin_AV_dout_mask
      );

    MPAR_L1D1EFGHin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1D1EFGHin_wea,
        addra     => MPAR_L1D1EFGHin_writeaddr,
        dina      => MPAR_L1D1EFGHin_din,
        wea_out       => MPAR_L1D1EFGHin_wea_delay,
        addra_out     => MPAR_L1D1EFGHin_writeaddr_delay,
        dina_out      => MPAR_L1D1EFGHin_din_delay,
        done       => PC_start,
        start      => MPAR_L1D1EFGHin_start
      );

    MPAR_L2D1ABCDin : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L2D1ABCDin"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L2D1ABCDin_wea_delay,
        addra     => MPAR_L2D1ABCDin_writeaddr_delay,
        dina      => MPAR_L2D1ABCDin_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L2D1ABCDin_V_readaddr,
        doutb     => MPAR_L2D1ABCDin_V_dout,
        sync_nent => MPAR_L2D1ABCDin_start,
        nent_o    => MPAR_L2D1ABCDin_AV_dout_nent,
        mask_o    => MPAR_L2D1ABCDin_AV_dout_mask
      );

    MPAR_L2D1ABCDin_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L2D1ABCDin_wea,
        addra     => MPAR_L2D1ABCDin_writeaddr,
        dina      => MPAR_L2D1ABCDin_din,
        wea_out       => MPAR_L2D1ABCDin_wea_delay,
        addra_out     => MPAR_L2D1ABCDin_writeaddr_delay,
        dina_out      => MPAR_L2D1ABCDin_din_delay,
        done       => PC_start,
        start      => MPAR_L2D1ABCDin_start
      );

    MPAR_L1L2ABC : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2ABC"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2ABC_wea_delay,
        addra     => MPAR_L1L2ABC_writeaddr_delay,
        dina      => MPAR_L1L2ABC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2ABC_V_readaddr,
        doutb     => MPAR_L1L2ABC_V_dout,
        sync_nent => MPAR_L1L2ABC_start,
        nent_o    => open
      );

    MPAR_L1L2ABC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2ABC_wea,
        addra     => MPAR_L1L2ABC_writeaddr,
        dina      => MPAR_L1L2ABC_din,
        wea_out       => MPAR_L1L2ABC_wea_delay,
        addra_out     => MPAR_L1L2ABC_writeaddr_delay,
        dina_out      => MPAR_L1L2ABC_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2ABC_start
      );

    MPAR_L1L2DE : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2DE"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2DE_wea_delay,
        addra     => MPAR_L1L2DE_writeaddr_delay,
        dina      => MPAR_L1L2DE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2DE_V_readaddr,
        doutb     => MPAR_L1L2DE_V_dout,
        sync_nent => MPAR_L1L2DE_start,
        nent_o    => open
      );

    MPAR_L1L2DE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2DE_wea,
        addra     => MPAR_L1L2DE_writeaddr,
        dina      => MPAR_L1L2DE_din,
        wea_out       => MPAR_L1L2DE_wea_delay,
        addra_out     => MPAR_L1L2DE_writeaddr_delay,
        dina_out      => MPAR_L1L2DE_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2DE_start
      );

    MPAR_L1L2F : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2F"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2F_wea_delay,
        addra     => MPAR_L1L2F_writeaddr_delay,
        dina      => MPAR_L1L2F_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2F_V_readaddr,
        doutb     => MPAR_L1L2F_V_dout,
        sync_nent => MPAR_L1L2F_start,
        nent_o    => open
      );

    MPAR_L1L2F_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2F_wea,
        addra     => MPAR_L1L2F_writeaddr,
        dina      => MPAR_L1L2F_din,
        wea_out       => MPAR_L1L2F_wea_delay,
        addra_out     => MPAR_L1L2F_writeaddr_delay,
        dina_out      => MPAR_L1L2F_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2F_start
      );

    MPAR_L1L2G : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2G"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2G_wea_delay,
        addra     => MPAR_L1L2G_writeaddr_delay,
        dina      => MPAR_L1L2G_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2G_V_readaddr,
        doutb     => MPAR_L1L2G_V_dout,
        sync_nent => MPAR_L1L2G_start,
        nent_o    => open
      );

    MPAR_L1L2G_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2G_wea,
        addra     => MPAR_L1L2G_writeaddr,
        dina      => MPAR_L1L2G_din,
        wea_out       => MPAR_L1L2G_wea_delay,
        addra_out     => MPAR_L1L2G_writeaddr_delay,
        dina_out      => MPAR_L1L2G_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2G_start
      );

    MPAR_L1L2HI : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2HI"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2HI_wea_delay,
        addra     => MPAR_L1L2HI_writeaddr_delay,
        dina      => MPAR_L1L2HI_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2HI_V_readaddr,
        doutb     => MPAR_L1L2HI_V_dout,
        sync_nent => MPAR_L1L2HI_start,
        nent_o    => open
      );

    MPAR_L1L2HI_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2HI_wea,
        addra     => MPAR_L1L2HI_writeaddr,
        dina      => MPAR_L1L2HI_din,
        wea_out       => MPAR_L1L2HI_wea_delay,
        addra_out     => MPAR_L1L2HI_writeaddr_delay,
        dina_out      => MPAR_L1L2HI_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2HI_start
      );

    MPAR_L1L2JKL : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1L2JKL"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1L2JKL_wea_delay,
        addra     => MPAR_L1L2JKL_writeaddr_delay,
        dina      => MPAR_L1L2JKL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1L2JKL_V_readaddr,
        doutb     => MPAR_L1L2JKL_V_dout,
        sync_nent => MPAR_L1L2JKL_start,
        nent_o    => open
      );

    MPAR_L1L2JKL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1L2JKL_wea,
        addra     => MPAR_L1L2JKL_writeaddr,
        dina      => MPAR_L1L2JKL_din,
        wea_out       => MPAR_L1L2JKL_wea_delay,
        addra_out     => MPAR_L1L2JKL_writeaddr_delay,
        dina_out      => MPAR_L1L2JKL_din_delay,
        done       => PC_done,
        start      => MPAR_L1L2JKL_start
      );

    MPAR_L2L3ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L2L3ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L2L3ABCD_wea_delay,
        addra     => MPAR_L2L3ABCD_writeaddr_delay,
        dina      => MPAR_L2L3ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L2L3ABCD_V_readaddr,
        doutb     => MPAR_L2L3ABCD_V_dout,
        sync_nent => MPAR_L2L3ABCD_start,
        nent_o    => open
      );

    MPAR_L2L3ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L2L3ABCD_wea,
        addra     => MPAR_L2L3ABCD_writeaddr,
        dina      => MPAR_L2L3ABCD_din,
        wea_out       => MPAR_L2L3ABCD_wea_delay,
        addra_out     => MPAR_L2L3ABCD_writeaddr_delay,
        dina_out      => MPAR_L2L3ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_L2L3ABCD_start
      );

    MPAR_L3L4AB : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L3L4AB"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L3L4AB_wea_delay,
        addra     => MPAR_L3L4AB_writeaddr_delay,
        dina      => MPAR_L3L4AB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L3L4AB_V_readaddr,
        doutb     => MPAR_L3L4AB_V_dout,
        sync_nent => MPAR_L3L4AB_start,
        nent_o    => open
      );

    MPAR_L3L4AB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L3L4AB_wea,
        addra     => MPAR_L3L4AB_writeaddr,
        dina      => MPAR_L3L4AB_din,
        wea_out       => MPAR_L3L4AB_wea_delay,
        addra_out     => MPAR_L3L4AB_writeaddr_delay,
        dina_out      => MPAR_L3L4AB_din_delay,
        done       => PC_done,
        start      => MPAR_L3L4AB_start
      );

    MPAR_L3L4CD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L3L4CD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L3L4CD_wea_delay,
        addra     => MPAR_L3L4CD_writeaddr_delay,
        dina      => MPAR_L3L4CD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L3L4CD_V_readaddr,
        doutb     => MPAR_L3L4CD_V_dout,
        sync_nent => MPAR_L3L4CD_start,
        nent_o    => open
      );

    MPAR_L3L4CD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L3L4CD_wea,
        addra     => MPAR_L3L4CD_writeaddr,
        dina      => MPAR_L3L4CD_din,
        wea_out       => MPAR_L3L4CD_wea_delay,
        addra_out     => MPAR_L3L4CD_writeaddr_delay,
        dina_out      => MPAR_L3L4CD_din_delay,
        done       => PC_done,
        start      => MPAR_L3L4CD_start
      );

    MPAR_L5L6ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L5L6ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L5L6ABCD_wea_delay,
        addra     => MPAR_L5L6ABCD_writeaddr_delay,
        dina      => MPAR_L5L6ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L5L6ABCD_V_readaddr,
        doutb     => MPAR_L5L6ABCD_V_dout,
        sync_nent => MPAR_L5L6ABCD_start,
        nent_o    => open
      );

    MPAR_L5L6ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L5L6ABCD_wea,
        addra     => MPAR_L5L6ABCD_writeaddr,
        dina      => MPAR_L5L6ABCD_din,
        wea_out       => MPAR_L5L6ABCD_wea_delay,
        addra_out     => MPAR_L5L6ABCD_writeaddr_delay,
        dina_out      => MPAR_L5L6ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_L5L6ABCD_start
      );

    MPAR_D1D2ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_D1D2ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_D1D2ABCD_wea_delay,
        addra     => MPAR_D1D2ABCD_writeaddr_delay,
        dina      => MPAR_D1D2ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_D1D2ABCD_V_readaddr,
        doutb     => MPAR_D1D2ABCD_V_dout,
        sync_nent => MPAR_D1D2ABCD_start,
        nent_o    => open
      );

    MPAR_D1D2ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_D1D2ABCD_wea,
        addra     => MPAR_D1D2ABCD_writeaddr,
        dina      => MPAR_D1D2ABCD_din,
        wea_out       => MPAR_D1D2ABCD_wea_delay,
        addra_out     => MPAR_D1D2ABCD_writeaddr_delay,
        dina_out      => MPAR_D1D2ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_D1D2ABCD_start
      );

    MPAR_D3D4ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_D3D4ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_D3D4ABCD_wea_delay,
        addra     => MPAR_D3D4ABCD_writeaddr_delay,
        dina      => MPAR_D3D4ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_D3D4ABCD_V_readaddr,
        doutb     => MPAR_D3D4ABCD_V_dout,
        sync_nent => MPAR_D3D4ABCD_start,
        nent_o    => open
      );

    MPAR_D3D4ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_D3D4ABCD_wea,
        addra     => MPAR_D3D4ABCD_writeaddr,
        dina      => MPAR_D3D4ABCD_din,
        wea_out       => MPAR_D3D4ABCD_wea_delay,
        addra_out     => MPAR_D3D4ABCD_writeaddr_delay,
        dina_out      => MPAR_D3D4ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_D3D4ABCD_start
      );

    MPAR_L1D1ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1D1ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1D1ABCD_wea_delay,
        addra     => MPAR_L1D1ABCD_writeaddr_delay,
        dina      => MPAR_L1D1ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1D1ABCD_V_readaddr,
        doutb     => MPAR_L1D1ABCD_V_dout,
        sync_nent => MPAR_L1D1ABCD_start,
        nent_o    => open
      );

    MPAR_L1D1ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1D1ABCD_wea,
        addra     => MPAR_L1D1ABCD_writeaddr,
        dina      => MPAR_L1D1ABCD_din,
        wea_out       => MPAR_L1D1ABCD_wea_delay,
        addra_out     => MPAR_L1D1ABCD_writeaddr_delay,
        dina_out      => MPAR_L1D1ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_L1D1ABCD_start
      );

    MPAR_L1D1EFGH : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L1D1EFGH"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L1D1EFGH_wea_delay,
        addra     => MPAR_L1D1EFGH_writeaddr_delay,
        dina      => MPAR_L1D1EFGH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L1D1EFGH_V_readaddr,
        doutb     => MPAR_L1D1EFGH_V_dout,
        sync_nent => MPAR_L1D1EFGH_start,
        nent_o    => open
      );

    MPAR_L1D1EFGH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L1D1EFGH_wea,
        addra     => MPAR_L1D1EFGH_writeaddr,
        dina      => MPAR_L1D1EFGH_din,
        wea_out       => MPAR_L1D1EFGH_wea_delay,
        addra_out     => MPAR_L1D1EFGH_writeaddr_delay,
        dina_out      => MPAR_L1D1EFGH_din_delay,
        done       => PC_done,
        start      => MPAR_L1D1EFGH_start
      );

    MPAR_L2D1ABCD : entity work.tf_mem_tpar
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPAR_L2D1ABCD"
      )
      port map (
        clka      => clk,
        wea       => MPAR_L2D1ABCD_wea_delay,
        addra     => MPAR_L2D1ABCD_writeaddr_delay,
        dina      => MPAR_L2D1ABCD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPAR_L2D1ABCD_V_readaddr,
        doutb     => MPAR_L2D1ABCD_V_dout,
        sync_nent => MPAR_L2D1ABCD_start,
        nent_o    => open
      );

    MPAR_L2D1ABCD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 32,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => MPAR_L2D1ABCD_wea,
        addra     => MPAR_L2D1ABCD_writeaddr,
        dina      => MPAR_L2D1ABCD_din,
        wea_out       => MPAR_L2D1ABCD_wea_delay,
        addra_out     => MPAR_L2D1ABCD_writeaddr_delay,
        dina_out      => MPAR_L2D1ABCD_din_delay,
        done       => PC_done,
        start      => MPAR_L2D1ABCD_start
      );

    MPROJ_L2L3ABCD_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIA_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIA_start
      );

    MPROJ_L3L4AB_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHIA_start,
        nent_o    => MPROJ_L3L4AB_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHIA_wea,
        addra     => MPROJ_L3L4AB_L1PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHIA_din,
        wea_out       => MPROJ_L3L4AB_L1PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHIA_start
      );

    MPROJ_L5L6ABCD_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIA_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIA_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIA_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIA_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIA_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIA_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIA_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIA_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIA_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIA_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIA_start
      );

    MPROJ_D1D2ABCD_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIA_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIA_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIA_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIA_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIA_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIA_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIA_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIA_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIA_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIA_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIA_start
      );

    MPROJ_D3D4ABCD_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIA_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIA_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIA_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIA_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIA_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIA_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIA_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIA_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIA_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIA_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIA_start
      );

    MPROJ_L2D1ABCD_L1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIA_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIA_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIA_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIA_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIA_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIA_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIA_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIA_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIA_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIA_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIA_start
      );

    MPROJ_L2L3ABCD_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIB_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIB_start
      );

    MPROJ_L3L4AB_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHIB_start,
        nent_o    => MPROJ_L3L4AB_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHIB_wea,
        addra     => MPROJ_L3L4AB_L1PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHIB_din,
        wea_out       => MPROJ_L3L4AB_L1PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHIB_start
      );

    MPROJ_L5L6ABCD_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIB_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIB_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIB_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIB_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIB_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIB_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIB_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIB_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIB_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIB_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIB_start
      );

    MPROJ_D1D2ABCD_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIB_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIB_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIB_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIB_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIB_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIB_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIB_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIB_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIB_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIB_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIB_start
      );

    MPROJ_D3D4ABCD_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIB_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIB_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIB_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIB_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIB_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIB_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIB_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIB_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIB_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIB_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIB_start
      );

    MPROJ_L2D1ABCD_L1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIB_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIB_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIB_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIB_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIB_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIB_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIB_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIB_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIB_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIB_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIB_start
      );

    MPROJ_L2L3ABCD_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIC_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIC_start
      );

    MPROJ_L3L4AB_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHIC_start,
        nent_o    => MPROJ_L3L4AB_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHIC_wea,
        addra     => MPROJ_L3L4AB_L1PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHIC_din,
        wea_out       => MPROJ_L3L4AB_L1PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHIC_start
      );

    MPROJ_L5L6ABCD_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIC_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIC_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIC_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIC_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIC_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIC_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIC_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIC_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIC_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIC_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIC_start
      );

    MPROJ_D1D2ABCD_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIC_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIC_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIC_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIC_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIC_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIC_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIC_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIC_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIC_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIC_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIC_start
      );

    MPROJ_D3D4ABCD_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIC_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIC_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIC_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIC_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIC_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIC_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIC_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIC_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIC_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIC_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIC_start
      );

    MPROJ_L2D1ABCD_L1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIC_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIC_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIC_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIC_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIC_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIC_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIC_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIC_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIC_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIC_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIC_start
      );

    MPROJ_L2L3ABCD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHID_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHID_wea,
        addra     => MPROJ_L2L3ABCD_L1PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHID_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHID_start
      );

    MPROJ_L3L4AB_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHID_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHID_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHID_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHID_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHID_start,
        nent_o    => MPROJ_L3L4AB_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHID_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHID_wea,
        addra     => MPROJ_L3L4AB_L1PHID_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHID_din,
        wea_out       => MPROJ_L3L4AB_L1PHID_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHID_start
      );

    MPROJ_L3L4CD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L1PHID_wea_delay,
        addra     => MPROJ_L3L4CD_L1PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L1PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_L1PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_L1PHID_start,
        nent_o    => MPROJ_L3L4CD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L1PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L1PHID_wea,
        addra     => MPROJ_L3L4CD_L1PHID_writeaddr,
        dina      => MPROJ_L3L4CD_L1PHID_din,
        wea_out       => MPROJ_L3L4CD_L1PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L1PHID_start
      );

    MPROJ_L5L6ABCD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHID_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHID_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHID_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHID_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHID_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHID_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHID_wea,
        addra     => MPROJ_L5L6ABCD_L1PHID_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHID_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHID_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHID_start
      );

    MPROJ_D1D2ABCD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHID_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHID_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHID_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHID_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHID_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHID_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHID_wea,
        addra     => MPROJ_D1D2ABCD_L1PHID_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHID_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHID_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHID_start
      );

    MPROJ_D3D4ABCD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHID_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHID_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHID_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHID_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHID_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHID_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHID_wea,
        addra     => MPROJ_D3D4ABCD_L1PHID_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHID_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHID_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHID_start
      );

    MPROJ_L2D1ABCD_L1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHID_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHID_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHID_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHID_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHID_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHID_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHID_wea,
        addra     => MPROJ_L2D1ABCD_L1PHID_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHID_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHID_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHID_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHID_start
      );

    MPROJ_L2L3ABCD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIE_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIE_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIE_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIE_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIE_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIE_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIE_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIE_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIE_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIE_start
      );

    MPROJ_L3L4AB_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHIE_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHIE_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHIE_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHIE_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHIE_start,
        nent_o    => MPROJ_L3L4AB_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHIE_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHIE_wea,
        addra     => MPROJ_L3L4AB_L1PHIE_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHIE_din,
        wea_out       => MPROJ_L3L4AB_L1PHIE_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHIE_start
      );

    MPROJ_L3L4CD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L1PHIE_wea_delay,
        addra     => MPROJ_L3L4CD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L1PHIE_V_readaddr,
        doutb     => MPROJ_L3L4CD_L1PHIE_V_dout,
        sync_nent => MPROJ_L3L4CD_L1PHIE_start,
        nent_o    => MPROJ_L3L4CD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L1PHIE_AV_dout_mask
      );

    MPROJ_L3L4CD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L1PHIE_wea,
        addra     => MPROJ_L3L4CD_L1PHIE_writeaddr,
        dina      => MPROJ_L3L4CD_L1PHIE_din,
        wea_out       => MPROJ_L3L4CD_L1PHIE_wea_delay,
        addra_out     => MPROJ_L3L4CD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L1PHIE_start
      );

    MPROJ_L5L6ABCD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIE_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIE_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIE_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIE_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIE_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIE_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIE_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIE_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIE_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIE_start
      );

    MPROJ_D1D2ABCD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIE_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIE_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIE_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIE_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIE_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIE_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIE_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIE_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIE_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIE_start
      );

    MPROJ_D3D4ABCD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIE_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIE_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIE_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIE_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIE_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIE_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIE_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIE_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIE_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIE_start
      );

    MPROJ_L2D1ABCD_L1PHIE : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIE_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIE_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIE_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIE_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIE_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIE_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIE_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIE_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIE_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIE_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIE_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIE_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIE_start
      );

    MPROJ_L2L3ABCD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIF_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIF_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIF_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIF_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIF_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIF_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIF_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIF_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIF_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIF_start
      );

    MPROJ_L3L4AB_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L1PHIF_wea_delay,
        addra     => MPROJ_L3L4AB_L1PHIF_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L1PHIF_V_readaddr,
        doutb     => MPROJ_L3L4AB_L1PHIF_V_dout,
        sync_nent => MPROJ_L3L4AB_L1PHIF_start,
        nent_o    => MPROJ_L3L4AB_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L1PHIF_AV_dout_mask
      );

    MPROJ_L3L4AB_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L1PHIF_wea,
        addra     => MPROJ_L3L4AB_L1PHIF_writeaddr,
        dina      => MPROJ_L3L4AB_L1PHIF_din,
        wea_out       => MPROJ_L3L4AB_L1PHIF_wea_delay,
        addra_out     => MPROJ_L3L4AB_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L1PHIF_start
      );

    MPROJ_L3L4CD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L1PHIF_wea_delay,
        addra     => MPROJ_L3L4CD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L1PHIF_V_readaddr,
        doutb     => MPROJ_L3L4CD_L1PHIF_V_dout,
        sync_nent => MPROJ_L3L4CD_L1PHIF_start,
        nent_o    => MPROJ_L3L4CD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L1PHIF_AV_dout_mask
      );

    MPROJ_L3L4CD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L1PHIF_wea,
        addra     => MPROJ_L3L4CD_L1PHIF_writeaddr,
        dina      => MPROJ_L3L4CD_L1PHIF_din,
        wea_out       => MPROJ_L3L4CD_L1PHIF_wea_delay,
        addra_out     => MPROJ_L3L4CD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L1PHIF_start
      );

    MPROJ_L5L6ABCD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIF_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIF_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIF_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIF_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIF_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIF_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIF_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIF_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIF_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIF_start
      );

    MPROJ_D1D2ABCD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIF_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIF_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIF_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIF_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIF_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIF_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIF_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIF_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIF_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIF_start
      );

    MPROJ_D3D4ABCD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIF_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIF_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIF_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIF_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIF_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIF_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIF_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIF_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIF_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIF_start
      );

    MPROJ_L2D1ABCD_L1PHIF : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIF_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIF_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIF_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIF_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIF_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIF_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIF_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIF_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIF_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIF_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIF_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIF_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIF_start
      );

    MPROJ_L2L3ABCD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIG_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIG_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIG_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIG_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIG_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIG_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIG_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIG_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIG_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIG_start
      );

    MPROJ_L3L4CD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L1PHIG_wea_delay,
        addra     => MPROJ_L3L4CD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L1PHIG_V_readaddr,
        doutb     => MPROJ_L3L4CD_L1PHIG_V_dout,
        sync_nent => MPROJ_L3L4CD_L1PHIG_start,
        nent_o    => MPROJ_L3L4CD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L1PHIG_AV_dout_mask
      );

    MPROJ_L3L4CD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L1PHIG_wea,
        addra     => MPROJ_L3L4CD_L1PHIG_writeaddr,
        dina      => MPROJ_L3L4CD_L1PHIG_din,
        wea_out       => MPROJ_L3L4CD_L1PHIG_wea_delay,
        addra_out     => MPROJ_L3L4CD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L1PHIG_start
      );

    MPROJ_L5L6ABCD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIG_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIG_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIG_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIG_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIG_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIG_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIG_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIG_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIG_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIG_start
      );

    MPROJ_D1D2ABCD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIG_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIG_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIG_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIG_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIG_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIG_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIG_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIG_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIG_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIG_start
      );

    MPROJ_D3D4ABCD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIG_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIG_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIG_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIG_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIG_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIG_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIG_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIG_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIG_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIG_start
      );

    MPROJ_L2D1ABCD_L1PHIG : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIG_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIG_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIG_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIG_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIG_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIG_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIG_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIG_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIG_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIG_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIG_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIG_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIG_start
      );

    MPROJ_L2L3ABCD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIH_wea_delay,
        addra     => MPROJ_L2L3ABCD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L1PHIH_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L1PHIH_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L1PHIH_start,
        nent_o    => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L1PHIH_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L1PHIH_wea,
        addra     => MPROJ_L2L3ABCD_L1PHIH_writeaddr,
        dina      => MPROJ_L2L3ABCD_L1PHIH_din,
        wea_out       => MPROJ_L2L3ABCD_L1PHIH_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L1PHIH_start
      );

    MPROJ_L3L4CD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L1PHIH_wea_delay,
        addra     => MPROJ_L3L4CD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L1PHIH_V_readaddr,
        doutb     => MPROJ_L3L4CD_L1PHIH_V_dout,
        sync_nent => MPROJ_L3L4CD_L1PHIH_start,
        nent_o    => MPROJ_L3L4CD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L1PHIH_AV_dout_mask
      );

    MPROJ_L3L4CD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L1PHIH_wea,
        addra     => MPROJ_L3L4CD_L1PHIH_writeaddr,
        dina      => MPROJ_L3L4CD_L1PHIH_din,
        wea_out       => MPROJ_L3L4CD_L1PHIH_wea_delay,
        addra_out     => MPROJ_L3L4CD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L1PHIH_start
      );

    MPROJ_L5L6ABCD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIH_wea_delay,
        addra     => MPROJ_L5L6ABCD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L1PHIH_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L1PHIH_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L1PHIH_start,
        nent_o    => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L1PHIH_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L1PHIH_wea,
        addra     => MPROJ_L5L6ABCD_L1PHIH_writeaddr,
        dina      => MPROJ_L5L6ABCD_L1PHIH_din,
        wea_out       => MPROJ_L5L6ABCD_L1PHIH_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L1PHIH_start
      );

    MPROJ_D1D2ABCD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIH_wea_delay,
        addra     => MPROJ_D1D2ABCD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L1PHIH_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L1PHIH_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L1PHIH_start,
        nent_o    => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L1PHIH_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L1PHIH_wea,
        addra     => MPROJ_D1D2ABCD_L1PHIH_writeaddr,
        dina      => MPROJ_D1D2ABCD_L1PHIH_din,
        wea_out       => MPROJ_D1D2ABCD_L1PHIH_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L1PHIH_start
      );

    MPROJ_D3D4ABCD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIH_wea_delay,
        addra     => MPROJ_D3D4ABCD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_L1PHIH_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_L1PHIH_V_dout,
        sync_nent => MPROJ_D3D4ABCD_L1PHIH_start,
        nent_o    => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_L1PHIH_AV_dout_mask
      );

    MPROJ_D3D4ABCD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_L1PHIH_wea,
        addra     => MPROJ_D3D4ABCD_L1PHIH_writeaddr,
        dina      => MPROJ_D3D4ABCD_L1PHIH_din,
        wea_out       => MPROJ_D3D4ABCD_L1PHIH_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_L1PHIH_start
      );

    MPROJ_L2D1ABCD_L1PHIH : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIH_wea_delay,
        addra     => MPROJ_L2D1ABCD_L1PHIH_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_L1PHIH_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_L1PHIH_V_dout,
        sync_nent => MPROJ_L2D1ABCD_L1PHIH_start,
        nent_o    => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_L1PHIH_AV_dout_mask
      );

    MPROJ_L2D1ABCD_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_L1PHIH_wea,
        addra     => MPROJ_L2D1ABCD_L1PHIH_writeaddr,
        dina      => MPROJ_L2D1ABCD_L1PHIH_din,
        wea_out       => MPROJ_L2D1ABCD_L1PHIH_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_L1PHIH_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_L1PHIH_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_L1PHIH_start
      );

    MPROJ_L3L4AB_L2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L2PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_L2PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L2PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_L2PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_L2PHIA_start,
        nent_o    => MPROJ_L3L4AB_L2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L2PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_L2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L2PHIA_wea,
        addra     => MPROJ_L3L4AB_L2PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_L2PHIA_din,
        wea_out       => MPROJ_L3L4AB_L2PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_L2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L2PHIA_start
      );

    MPROJ_L5L6ABCD_L2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIA_wea_delay,
        addra     => MPROJ_L5L6ABCD_L2PHIA_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L2PHIA_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L2PHIA_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L2PHIA_start,
        nent_o    => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L2PHIA_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIA_wea,
        addra     => MPROJ_L5L6ABCD_L2PHIA_writeaddr,
        dina      => MPROJ_L5L6ABCD_L2PHIA_din,
        wea_out       => MPROJ_L5L6ABCD_L2PHIA_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L2PHIA_start
      );

    MPROJ_D1D2ABCD_L2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIA_wea_delay,
        addra     => MPROJ_D1D2ABCD_L2PHIA_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L2PHIA_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L2PHIA_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L2PHIA_start,
        nent_o    => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L2PHIA_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIA_wea,
        addra     => MPROJ_D1D2ABCD_L2PHIA_writeaddr,
        dina      => MPROJ_D1D2ABCD_L2PHIA_din,
        wea_out       => MPROJ_D1D2ABCD_L2PHIA_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L2PHIA_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L2PHIA_start
      );

    MPROJ_L3L4AB_L2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L2PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_L2PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L2PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_L2PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_L2PHIB_start,
        nent_o    => MPROJ_L3L4AB_L2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L2PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L2PHIB_wea,
        addra     => MPROJ_L3L4AB_L2PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_L2PHIB_din,
        wea_out       => MPROJ_L3L4AB_L2PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_L2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L2PHIB_start
      );

    MPROJ_L3L4CD_L2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L2PHIB_wea_delay,
        addra     => MPROJ_L3L4CD_L2PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L2PHIB_V_readaddr,
        doutb     => MPROJ_L3L4CD_L2PHIB_V_dout,
        sync_nent => MPROJ_L3L4CD_L2PHIB_start,
        nent_o    => MPROJ_L3L4CD_L2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L2PHIB_AV_dout_mask
      );

    MPROJ_L3L4CD_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L2PHIB_wea,
        addra     => MPROJ_L3L4CD_L2PHIB_writeaddr,
        dina      => MPROJ_L3L4CD_L2PHIB_din,
        wea_out       => MPROJ_L3L4CD_L2PHIB_wea_delay,
        addra_out     => MPROJ_L3L4CD_L2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L2PHIB_start
      );

    MPROJ_L5L6ABCD_L2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIB_wea_delay,
        addra     => MPROJ_L5L6ABCD_L2PHIB_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L2PHIB_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L2PHIB_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L2PHIB_start,
        nent_o    => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L2PHIB_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIB_wea,
        addra     => MPROJ_L5L6ABCD_L2PHIB_writeaddr,
        dina      => MPROJ_L5L6ABCD_L2PHIB_din,
        wea_out       => MPROJ_L5L6ABCD_L2PHIB_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L2PHIB_start
      );

    MPROJ_D1D2ABCD_L2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIB_wea_delay,
        addra     => MPROJ_D1D2ABCD_L2PHIB_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L2PHIB_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L2PHIB_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L2PHIB_start,
        nent_o    => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L2PHIB_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIB_wea,
        addra     => MPROJ_D1D2ABCD_L2PHIB_writeaddr,
        dina      => MPROJ_D1D2ABCD_L2PHIB_din,
        wea_out       => MPROJ_D1D2ABCD_L2PHIB_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L2PHIB_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L2PHIB_start
      );

    MPROJ_L3L4AB_L2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L2PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_L2PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L2PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_L2PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_L2PHIC_start,
        nent_o    => MPROJ_L3L4AB_L2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L2PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L2PHIC_wea,
        addra     => MPROJ_L3L4AB_L2PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_L2PHIC_din,
        wea_out       => MPROJ_L3L4AB_L2PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_L2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L2PHIC_start
      );

    MPROJ_L3L4CD_L2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L2PHIC_wea_delay,
        addra     => MPROJ_L3L4CD_L2PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L2PHIC_V_readaddr,
        doutb     => MPROJ_L3L4CD_L2PHIC_V_dout,
        sync_nent => MPROJ_L3L4CD_L2PHIC_start,
        nent_o    => MPROJ_L3L4CD_L2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L2PHIC_AV_dout_mask
      );

    MPROJ_L3L4CD_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L2PHIC_wea,
        addra     => MPROJ_L3L4CD_L2PHIC_writeaddr,
        dina      => MPROJ_L3L4CD_L2PHIC_din,
        wea_out       => MPROJ_L3L4CD_L2PHIC_wea_delay,
        addra_out     => MPROJ_L3L4CD_L2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L2PHIC_start
      );

    MPROJ_L5L6ABCD_L2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIC_wea_delay,
        addra     => MPROJ_L5L6ABCD_L2PHIC_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L2PHIC_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L2PHIC_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L2PHIC_start,
        nent_o    => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L2PHIC_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHIC_wea,
        addra     => MPROJ_L5L6ABCD_L2PHIC_writeaddr,
        dina      => MPROJ_L5L6ABCD_L2PHIC_din,
        wea_out       => MPROJ_L5L6ABCD_L2PHIC_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L2PHIC_start
      );

    MPROJ_D1D2ABCD_L2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIC_wea_delay,
        addra     => MPROJ_D1D2ABCD_L2PHIC_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L2PHIC_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L2PHIC_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L2PHIC_start,
        nent_o    => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L2PHIC_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHIC_wea,
        addra     => MPROJ_D1D2ABCD_L2PHIC_writeaddr,
        dina      => MPROJ_D1D2ABCD_L2PHIC_din,
        wea_out       => MPROJ_D1D2ABCD_L2PHIC_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L2PHIC_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L2PHIC_start
      );

    MPROJ_L3L4CD_L2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L2PHID_wea_delay,
        addra     => MPROJ_L3L4CD_L2PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L2PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_L2PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_L2PHID_start,
        nent_o    => MPROJ_L3L4CD_L2PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L2PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_L2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L2PHID_wea,
        addra     => MPROJ_L3L4CD_L2PHID_writeaddr,
        dina      => MPROJ_L3L4CD_L2PHID_din,
        wea_out       => MPROJ_L3L4CD_L2PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_L2PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L2PHID_start
      );

    MPROJ_L5L6ABCD_L2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHID_wea_delay,
        addra     => MPROJ_L5L6ABCD_L2PHID_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L2PHID_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L2PHID_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L2PHID_start,
        nent_o    => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L2PHID_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L2PHID_wea,
        addra     => MPROJ_L5L6ABCD_L2PHID_writeaddr,
        dina      => MPROJ_L5L6ABCD_L2PHID_din,
        wea_out       => MPROJ_L5L6ABCD_L2PHID_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L2PHID_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L2PHID_start
      );

    MPROJ_D1D2ABCD_L2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_L2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHID_wea_delay,
        addra     => MPROJ_D1D2ABCD_L2PHID_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_L2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_L2PHID_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_L2PHID_V_dout,
        sync_nent => MPROJ_D1D2ABCD_L2PHID_start,
        nent_o    => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_L2PHID_AV_dout_mask
      );

    MPROJ_D1D2ABCD_L2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_L2PHID_wea,
        addra     => MPROJ_D1D2ABCD_L2PHID_writeaddr,
        dina      => MPROJ_D1D2ABCD_L2PHID_din,
        wea_out       => MPROJ_D1D2ABCD_L2PHID_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_L2PHID_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_L2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_L2PHID_start
      );

    MPROJ_L1L2ABC_L3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L3PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_L3PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L3PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L3PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_L3PHIA_start,
        nent_o    => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L3PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_L3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L3PHIA_wea,
        addra     => MPROJ_L1L2ABC_L3PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_L3PHIA_din,
        wea_out       => MPROJ_L1L2ABC_L3PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L3PHIA_start
      );

    MPROJ_L1L2DE_L3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L3PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_L3PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L3PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_L3PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_L3PHIA_start,
        nent_o    => MPROJ_L1L2DE_L3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L3PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_L3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L3PHIA_wea,
        addra     => MPROJ_L1L2DE_L3PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_L3PHIA_din,
        wea_out       => MPROJ_L1L2DE_L3PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_L3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L3PHIA_start
      );

    MPROJ_L5L6ABCD_L3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIA_wea_delay,
        addra     => MPROJ_L5L6ABCD_L3PHIA_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L3PHIA_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L3PHIA_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L3PHIA_start,
        nent_o    => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L3PHIA_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIA_wea,
        addra     => MPROJ_L5L6ABCD_L3PHIA_writeaddr,
        dina      => MPROJ_L5L6ABCD_L3PHIA_din,
        wea_out       => MPROJ_L5L6ABCD_L3PHIA_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L3PHIA_start
      );

    MPROJ_L1L2ABC_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L3PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L3PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_L3PHIB_start,
        nent_o    => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L3PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L3PHIB_wea,
        addra     => MPROJ_L1L2ABC_L3PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_L3PHIB_din,
        wea_out       => MPROJ_L1L2ABC_L3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L3PHIB_start
      );

    MPROJ_L1L2DE_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L3PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_L3PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_L3PHIB_start,
        nent_o    => MPROJ_L1L2DE_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L3PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L3PHIB_wea,
        addra     => MPROJ_L1L2DE_L3PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_L3PHIB_din,
        wea_out       => MPROJ_L1L2DE_L3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L3PHIB_start
      );

    MPROJ_L1L2F_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L3PHIB_wea_delay,
        addra     => MPROJ_L1L2F_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_L3PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_L3PHIB_start,
        nent_o    => MPROJ_L1L2F_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L3PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L3PHIB_wea,
        addra     => MPROJ_L1L2F_L3PHIB_writeaddr,
        dina      => MPROJ_L1L2F_L3PHIB_din,
        wea_out       => MPROJ_L1L2F_L3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L3PHIB_start
      );

    MPROJ_L1L2G_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L3PHIB_wea_delay,
        addra     => MPROJ_L1L2G_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_L3PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_L3PHIB_start,
        nent_o    => MPROJ_L1L2G_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L3PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L3PHIB_wea,
        addra     => MPROJ_L1L2G_L3PHIB_writeaddr,
        dina      => MPROJ_L1L2G_L3PHIB_din,
        wea_out       => MPROJ_L1L2G_L3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L3PHIB_start
      );

    MPROJ_L1L2HI_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L3PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_L3PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_L3PHIB_start,
        nent_o    => MPROJ_L1L2HI_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L3PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L3PHIB_wea,
        addra     => MPROJ_L1L2HI_L3PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_L3PHIB_din,
        wea_out       => MPROJ_L1L2HI_L3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L3PHIB_start
      );

    MPROJ_L5L6ABCD_L3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIB_wea_delay,
        addra     => MPROJ_L5L6ABCD_L3PHIB_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L3PHIB_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L3PHIB_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L3PHIB_start,
        nent_o    => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L3PHIB_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIB_wea,
        addra     => MPROJ_L5L6ABCD_L3PHIB_writeaddr,
        dina      => MPROJ_L5L6ABCD_L3PHIB_din,
        wea_out       => MPROJ_L5L6ABCD_L3PHIB_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L3PHIB_start
      );

    MPROJ_L1L2DE_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L3PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_L3PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_L3PHIC_start,
        nent_o    => MPROJ_L1L2DE_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L3PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L3PHIC_wea,
        addra     => MPROJ_L1L2DE_L3PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_L3PHIC_din,
        wea_out       => MPROJ_L1L2DE_L3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L3PHIC_start
      );

    MPROJ_L1L2F_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L3PHIC_wea_delay,
        addra     => MPROJ_L1L2F_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_L3PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_L3PHIC_start,
        nent_o    => MPROJ_L1L2F_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L3PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L3PHIC_wea,
        addra     => MPROJ_L1L2F_L3PHIC_writeaddr,
        dina      => MPROJ_L1L2F_L3PHIC_din,
        wea_out       => MPROJ_L1L2F_L3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L3PHIC_start
      );

    MPROJ_L1L2G_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L3PHIC_wea_delay,
        addra     => MPROJ_L1L2G_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_L3PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_L3PHIC_start,
        nent_o    => MPROJ_L1L2G_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L3PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L3PHIC_wea,
        addra     => MPROJ_L1L2G_L3PHIC_writeaddr,
        dina      => MPROJ_L1L2G_L3PHIC_din,
        wea_out       => MPROJ_L1L2G_L3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L3PHIC_start
      );

    MPROJ_L1L2HI_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L3PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_L3PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_L3PHIC_start,
        nent_o    => MPROJ_L1L2HI_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L3PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L3PHIC_wea,
        addra     => MPROJ_L1L2HI_L3PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_L3PHIC_din,
        wea_out       => MPROJ_L1L2HI_L3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L3PHIC_start
      );

    MPROJ_L1L2JKL_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L3PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L3PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_L3PHIC_start,
        nent_o    => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L3PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L3PHIC_wea,
        addra     => MPROJ_L1L2JKL_L3PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_L3PHIC_din,
        wea_out       => MPROJ_L1L2JKL_L3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L3PHIC_start
      );

    MPROJ_L5L6ABCD_L3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIC_wea_delay,
        addra     => MPROJ_L5L6ABCD_L3PHIC_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L3PHIC_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L3PHIC_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L3PHIC_start,
        nent_o    => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L3PHIC_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHIC_wea,
        addra     => MPROJ_L5L6ABCD_L3PHIC_writeaddr,
        dina      => MPROJ_L5L6ABCD_L3PHIC_din,
        wea_out       => MPROJ_L5L6ABCD_L3PHIC_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L3PHIC_start
      );

    MPROJ_L1L2HI_L3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L3PHID_wea_delay,
        addra     => MPROJ_L1L2HI_L3PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L3PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_L3PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_L3PHID_start,
        nent_o    => MPROJ_L1L2HI_L3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L3PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_L3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L3PHID_wea,
        addra     => MPROJ_L1L2HI_L3PHID_writeaddr,
        dina      => MPROJ_L1L2HI_L3PHID_din,
        wea_out       => MPROJ_L1L2HI_L3PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_L3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L3PHID_start
      );

    MPROJ_L1L2JKL_L3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L3PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_L3PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L3PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L3PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_L3PHID_start,
        nent_o    => MPROJ_L1L2JKL_L3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L3PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_L3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L3PHID_wea,
        addra     => MPROJ_L1L2JKL_L3PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_L3PHID_din,
        wea_out       => MPROJ_L1L2JKL_L3PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L3PHID_start
      );

    MPROJ_L5L6ABCD_L3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHID_wea_delay,
        addra     => MPROJ_L5L6ABCD_L3PHID_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L3PHID_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L3PHID_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L3PHID_start,
        nent_o    => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L3PHID_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 60
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L3PHID_wea,
        addra     => MPROJ_L5L6ABCD_L3PHID_writeaddr,
        dina      => MPROJ_L5L6ABCD_L3PHID_din,
        wea_out       => MPROJ_L5L6ABCD_L3PHID_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L3PHID_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L3PHID_start
      );

    MPROJ_L1L2ABC_L4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L4PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_L4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L4PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_L4PHIA_start,
        nent_o    => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L4PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L4PHIA_wea,
        addra     => MPROJ_L1L2ABC_L4PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_L4PHIA_din,
        wea_out       => MPROJ_L1L2ABC_L4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L4PHIA_start
      );

    MPROJ_L1L2DE_L4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L4PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_L4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_L4PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_L4PHIA_start,
        nent_o    => MPROJ_L1L2DE_L4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L4PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L4PHIA_wea,
        addra     => MPROJ_L1L2DE_L4PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_L4PHIA_din,
        wea_out       => MPROJ_L1L2DE_L4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_L4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L4PHIA_start
      );

    MPROJ_L1L2F_L4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L4PHIA_wea_delay,
        addra     => MPROJ_L1L2F_L4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_L4PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_L4PHIA_start,
        nent_o    => MPROJ_L1L2F_L4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L4PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L4PHIA_wea,
        addra     => MPROJ_L1L2F_L4PHIA_writeaddr,
        dina      => MPROJ_L1L2F_L4PHIA_din,
        wea_out       => MPROJ_L1L2F_L4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_L4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L4PHIA_start
      );

    MPROJ_L2L3ABCD_L4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_L4PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L4PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L4PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L4PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L4PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIA_wea,
        addra     => MPROJ_L2L3ABCD_L4PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_L4PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_L4PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L4PHIA_start
      );

    MPROJ_L5L6ABCD_L4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIA_wea_delay,
        addra     => MPROJ_L5L6ABCD_L4PHIA_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L4PHIA_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L4PHIA_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L4PHIA_start,
        nent_o    => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L4PHIA_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIA_wea,
        addra     => MPROJ_L5L6ABCD_L4PHIA_writeaddr,
        dina      => MPROJ_L5L6ABCD_L4PHIA_din,
        wea_out       => MPROJ_L5L6ABCD_L4PHIA_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L4PHIA_start
      );

    MPROJ_L1L2ABC_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L4PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L4PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_L4PHIB_start,
        nent_o    => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L4PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L4PHIB_wea,
        addra     => MPROJ_L1L2ABC_L4PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_L4PHIB_din,
        wea_out       => MPROJ_L1L2ABC_L4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L4PHIB_start
      );

    MPROJ_L1L2DE_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L4PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_L4PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_L4PHIB_start,
        nent_o    => MPROJ_L1L2DE_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L4PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L4PHIB_wea,
        addra     => MPROJ_L1L2DE_L4PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_L4PHIB_din,
        wea_out       => MPROJ_L1L2DE_L4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L4PHIB_start
      );

    MPROJ_L1L2F_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L4PHIB_wea_delay,
        addra     => MPROJ_L1L2F_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_L4PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_L4PHIB_start,
        nent_o    => MPROJ_L1L2F_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L4PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L4PHIB_wea,
        addra     => MPROJ_L1L2F_L4PHIB_writeaddr,
        dina      => MPROJ_L1L2F_L4PHIB_din,
        wea_out       => MPROJ_L1L2F_L4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L4PHIB_start
      );

    MPROJ_L1L2G_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L4PHIB_wea_delay,
        addra     => MPROJ_L1L2G_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_L4PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_L4PHIB_start,
        nent_o    => MPROJ_L1L2G_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L4PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L4PHIB_wea,
        addra     => MPROJ_L1L2G_L4PHIB_writeaddr,
        dina      => MPROJ_L1L2G_L4PHIB_din,
        wea_out       => MPROJ_L1L2G_L4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L4PHIB_start
      );

    MPROJ_L1L2HI_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L4PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_L4PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_L4PHIB_start,
        nent_o    => MPROJ_L1L2HI_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L4PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L4PHIB_wea,
        addra     => MPROJ_L1L2HI_L4PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_L4PHIB_din,
        wea_out       => MPROJ_L1L2HI_L4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L4PHIB_start
      );

    MPROJ_L2L3ABCD_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L4PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L4PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L4PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L4PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIB_wea,
        addra     => MPROJ_L2L3ABCD_L4PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_L4PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_L4PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L4PHIB_start
      );

    MPROJ_L5L6ABCD_L4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIB_wea_delay,
        addra     => MPROJ_L5L6ABCD_L4PHIB_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L4PHIB_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L4PHIB_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L4PHIB_start,
        nent_o    => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L4PHIB_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIB_wea,
        addra     => MPROJ_L5L6ABCD_L4PHIB_writeaddr,
        dina      => MPROJ_L5L6ABCD_L4PHIB_din,
        wea_out       => MPROJ_L5L6ABCD_L4PHIB_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L4PHIB_start
      );

    MPROJ_L1L2DE_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L4PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_L4PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_L4PHIC_start,
        nent_o    => MPROJ_L1L2DE_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L4PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L4PHIC_wea,
        addra     => MPROJ_L1L2DE_L4PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_L4PHIC_din,
        wea_out       => MPROJ_L1L2DE_L4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L4PHIC_start
      );

    MPROJ_L1L2F_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L4PHIC_wea_delay,
        addra     => MPROJ_L1L2F_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_L4PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_L4PHIC_start,
        nent_o    => MPROJ_L1L2F_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L4PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L4PHIC_wea,
        addra     => MPROJ_L1L2F_L4PHIC_writeaddr,
        dina      => MPROJ_L1L2F_L4PHIC_din,
        wea_out       => MPROJ_L1L2F_L4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L4PHIC_start
      );

    MPROJ_L1L2G_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L4PHIC_wea_delay,
        addra     => MPROJ_L1L2G_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_L4PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_L4PHIC_start,
        nent_o    => MPROJ_L1L2G_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L4PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L4PHIC_wea,
        addra     => MPROJ_L1L2G_L4PHIC_writeaddr,
        dina      => MPROJ_L1L2G_L4PHIC_din,
        wea_out       => MPROJ_L1L2G_L4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L4PHIC_start
      );

    MPROJ_L1L2HI_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L4PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_L4PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_L4PHIC_start,
        nent_o    => MPROJ_L1L2HI_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L4PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L4PHIC_wea,
        addra     => MPROJ_L1L2HI_L4PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_L4PHIC_din,
        wea_out       => MPROJ_L1L2HI_L4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L4PHIC_start
      );

    MPROJ_L1L2JKL_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L4PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L4PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_L4PHIC_start,
        nent_o    => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L4PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L4PHIC_wea,
        addra     => MPROJ_L1L2JKL_L4PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_L4PHIC_din,
        wea_out       => MPROJ_L1L2JKL_L4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L4PHIC_start
      );

    MPROJ_L2L3ABCD_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L4PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L4PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L4PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L4PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHIC_wea,
        addra     => MPROJ_L2L3ABCD_L4PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_L4PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_L4PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L4PHIC_start
      );

    MPROJ_L5L6ABCD_L4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIC_wea_delay,
        addra     => MPROJ_L5L6ABCD_L4PHIC_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L4PHIC_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L4PHIC_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L4PHIC_start,
        nent_o    => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L4PHIC_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHIC_wea,
        addra     => MPROJ_L5L6ABCD_L4PHIC_writeaddr,
        dina      => MPROJ_L5L6ABCD_L4PHIC_din,
        wea_out       => MPROJ_L5L6ABCD_L4PHIC_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L4PHIC_start
      );

    MPROJ_L1L2G_L4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L4PHID_wea_delay,
        addra     => MPROJ_L1L2G_L4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L4PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_L4PHID_V_dout,
        sync_nent => MPROJ_L1L2G_L4PHID_start,
        nent_o    => MPROJ_L1L2G_L4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L4PHID_AV_dout_mask
      );

    MPROJ_L1L2G_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L4PHID_wea,
        addra     => MPROJ_L1L2G_L4PHID_writeaddr,
        dina      => MPROJ_L1L2G_L4PHID_din,
        wea_out       => MPROJ_L1L2G_L4PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_L4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L4PHID_start
      );

    MPROJ_L1L2HI_L4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L4PHID_wea_delay,
        addra     => MPROJ_L1L2HI_L4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L4PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_L4PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_L4PHID_start,
        nent_o    => MPROJ_L1L2HI_L4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L4PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L4PHID_wea,
        addra     => MPROJ_L1L2HI_L4PHID_writeaddr,
        dina      => MPROJ_L1L2HI_L4PHID_din,
        wea_out       => MPROJ_L1L2HI_L4PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_L4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L4PHID_start
      );

    MPROJ_L1L2JKL_L4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L4PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_L4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L4PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L4PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_L4PHID_start,
        nent_o    => MPROJ_L1L2JKL_L4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L4PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L4PHID_wea,
        addra     => MPROJ_L1L2JKL_L4PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_L4PHID_din,
        wea_out       => MPROJ_L1L2JKL_L4PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L4PHID_start
      );

    MPROJ_L2L3ABCD_L4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_L4PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L4PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L4PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L4PHID_start,
        nent_o    => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L4PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L4PHID_wea,
        addra     => MPROJ_L2L3ABCD_L4PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_L4PHID_din,
        wea_out       => MPROJ_L2L3ABCD_L4PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L4PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L4PHID_start
      );

    MPROJ_L5L6ABCD_L4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L5L6ABCD_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHID_wea_delay,
        addra     => MPROJ_L5L6ABCD_L4PHID_writeaddr_delay,
        dina      => MPROJ_L5L6ABCD_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L5L6ABCD_L4PHID_V_readaddr,
        doutb     => MPROJ_L5L6ABCD_L4PHID_V_dout,
        sync_nent => MPROJ_L5L6ABCD_L4PHID_start,
        nent_o    => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent,
        mask_o    => MPROJ_L5L6ABCD_L4PHID_AV_dout_mask
      );

    MPROJ_L5L6ABCD_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L5L6ABCD_L4PHID_wea,
        addra     => MPROJ_L5L6ABCD_L4PHID_writeaddr,
        dina      => MPROJ_L5L6ABCD_L4PHID_din,
        wea_out       => MPROJ_L5L6ABCD_L4PHID_wea_delay,
        addra_out     => MPROJ_L5L6ABCD_L4PHID_writeaddr_delay,
        dina_out      => MPROJ_L5L6ABCD_L4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L5L6ABCD_L4PHID_start
      );

    MPROJ_L1L2ABC_L5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L5PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_L5PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L5PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L5PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_L5PHIA_start,
        nent_o    => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L5PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L5PHIA_wea,
        addra     => MPROJ_L1L2ABC_L5PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_L5PHIA_din,
        wea_out       => MPROJ_L1L2ABC_L5PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L5PHIA_start
      );

    MPROJ_L1L2DE_L5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L5PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_L5PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L5PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_L5PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_L5PHIA_start,
        nent_o    => MPROJ_L1L2DE_L5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L5PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L5PHIA_wea,
        addra     => MPROJ_L1L2DE_L5PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_L5PHIA_din,
        wea_out       => MPROJ_L1L2DE_L5PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_L5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L5PHIA_start
      );

    MPROJ_L1L2F_L5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L5PHIA_wea_delay,
        addra     => MPROJ_L1L2F_L5PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L5PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_L5PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_L5PHIA_start,
        nent_o    => MPROJ_L1L2F_L5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L5PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L5PHIA_wea,
        addra     => MPROJ_L1L2F_L5PHIA_writeaddr,
        dina      => MPROJ_L1L2F_L5PHIA_din,
        wea_out       => MPROJ_L1L2F_L5PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_L5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L5PHIA_start
      );

    MPROJ_L2L3ABCD_L5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_L5PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L5PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L5PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L5PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L5PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIA_wea,
        addra     => MPROJ_L2L3ABCD_L5PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_L5PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_L5PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L5PHIA_start
      );

    MPROJ_L3L4AB_L5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L5PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_L5PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L5PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_L5PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_L5PHIA_start,
        nent_o    => MPROJ_L3L4AB_L5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L5PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L5PHIA_wea,
        addra     => MPROJ_L3L4AB_L5PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_L5PHIA_din,
        wea_out       => MPROJ_L3L4AB_L5PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_L5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L5PHIA_start
      );

    MPROJ_L1L2ABC_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L5PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L5PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L5PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_L5PHIB_start,
        nent_o    => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L5PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L5PHIB_wea,
        addra     => MPROJ_L1L2ABC_L5PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_L5PHIB_din,
        wea_out       => MPROJ_L1L2ABC_L5PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L5PHIB_start
      );

    MPROJ_L1L2DE_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L5PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L5PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_L5PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_L5PHIB_start,
        nent_o    => MPROJ_L1L2DE_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L5PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L5PHIB_wea,
        addra     => MPROJ_L1L2DE_L5PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_L5PHIB_din,
        wea_out       => MPROJ_L1L2DE_L5PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L5PHIB_start
      );

    MPROJ_L1L2F_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L5PHIB_wea_delay,
        addra     => MPROJ_L1L2F_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L5PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_L5PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_L5PHIB_start,
        nent_o    => MPROJ_L1L2F_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L5PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L5PHIB_wea,
        addra     => MPROJ_L1L2F_L5PHIB_writeaddr,
        dina      => MPROJ_L1L2F_L5PHIB_din,
        wea_out       => MPROJ_L1L2F_L5PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L5PHIB_start
      );

    MPROJ_L1L2G_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L5PHIB_wea_delay,
        addra     => MPROJ_L1L2G_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L5PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_L5PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_L5PHIB_start,
        nent_o    => MPROJ_L1L2G_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L5PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L5PHIB_wea,
        addra     => MPROJ_L1L2G_L5PHIB_writeaddr,
        dina      => MPROJ_L1L2G_L5PHIB_din,
        wea_out       => MPROJ_L1L2G_L5PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L5PHIB_start
      );

    MPROJ_L1L2HI_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L5PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L5PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_L5PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_L5PHIB_start,
        nent_o    => MPROJ_L1L2HI_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L5PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L5PHIB_wea,
        addra     => MPROJ_L1L2HI_L5PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_L5PHIB_din,
        wea_out       => MPROJ_L1L2HI_L5PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L5PHIB_start
      );

    MPROJ_L2L3ABCD_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L5PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L5PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L5PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L5PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIB_wea,
        addra     => MPROJ_L2L3ABCD_L5PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_L5PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_L5PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L5PHIB_start
      );

    MPROJ_L3L4AB_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L5PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L5PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_L5PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_L5PHIB_start,
        nent_o    => MPROJ_L3L4AB_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L5PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L5PHIB_wea,
        addra     => MPROJ_L3L4AB_L5PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_L5PHIB_din,
        wea_out       => MPROJ_L3L4AB_L5PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L5PHIB_start
      );

    MPROJ_L3L4CD_L5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L5PHIB_wea_delay,
        addra     => MPROJ_L3L4CD_L5PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L5PHIB_V_readaddr,
        doutb     => MPROJ_L3L4CD_L5PHIB_V_dout,
        sync_nent => MPROJ_L3L4CD_L5PHIB_start,
        nent_o    => MPROJ_L3L4CD_L5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L5PHIB_AV_dout_mask
      );

    MPROJ_L3L4CD_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L5PHIB_wea,
        addra     => MPROJ_L3L4CD_L5PHIB_writeaddr,
        dina      => MPROJ_L3L4CD_L5PHIB_din,
        wea_out       => MPROJ_L3L4CD_L5PHIB_wea_delay,
        addra_out     => MPROJ_L3L4CD_L5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L5PHIB_start
      );

    MPROJ_L1L2DE_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L5PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L5PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_L5PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_L5PHIC_start,
        nent_o    => MPROJ_L1L2DE_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L5PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L5PHIC_wea,
        addra     => MPROJ_L1L2DE_L5PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_L5PHIC_din,
        wea_out       => MPROJ_L1L2DE_L5PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L5PHIC_start
      );

    MPROJ_L1L2F_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L5PHIC_wea_delay,
        addra     => MPROJ_L1L2F_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L5PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_L5PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_L5PHIC_start,
        nent_o    => MPROJ_L1L2F_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L5PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L5PHIC_wea,
        addra     => MPROJ_L1L2F_L5PHIC_writeaddr,
        dina      => MPROJ_L1L2F_L5PHIC_din,
        wea_out       => MPROJ_L1L2F_L5PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L5PHIC_start
      );

    MPROJ_L1L2G_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L5PHIC_wea_delay,
        addra     => MPROJ_L1L2G_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L5PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_L5PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_L5PHIC_start,
        nent_o    => MPROJ_L1L2G_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L5PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L5PHIC_wea,
        addra     => MPROJ_L1L2G_L5PHIC_writeaddr,
        dina      => MPROJ_L1L2G_L5PHIC_din,
        wea_out       => MPROJ_L1L2G_L5PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L5PHIC_start
      );

    MPROJ_L1L2HI_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L5PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L5PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_L5PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_L5PHIC_start,
        nent_o    => MPROJ_L1L2HI_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L5PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L5PHIC_wea,
        addra     => MPROJ_L1L2HI_L5PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_L5PHIC_din,
        wea_out       => MPROJ_L1L2HI_L5PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L5PHIC_start
      );

    MPROJ_L1L2JKL_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L5PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L5PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L5PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_L5PHIC_start,
        nent_o    => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L5PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L5PHIC_wea,
        addra     => MPROJ_L1L2JKL_L5PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_L5PHIC_din,
        wea_out       => MPROJ_L1L2JKL_L5PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L5PHIC_start
      );

    MPROJ_L2L3ABCD_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L5PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L5PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L5PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L5PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHIC_wea,
        addra     => MPROJ_L2L3ABCD_L5PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_L5PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_L5PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L5PHIC_start
      );

    MPROJ_L3L4AB_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L5PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L5PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_L5PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_L5PHIC_start,
        nent_o    => MPROJ_L3L4AB_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L5PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L5PHIC_wea,
        addra     => MPROJ_L3L4AB_L5PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_L5PHIC_din,
        wea_out       => MPROJ_L3L4AB_L5PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L5PHIC_start
      );

    MPROJ_L3L4CD_L5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L5PHIC_wea_delay,
        addra     => MPROJ_L3L4CD_L5PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L5PHIC_V_readaddr,
        doutb     => MPROJ_L3L4CD_L5PHIC_V_dout,
        sync_nent => MPROJ_L3L4CD_L5PHIC_start,
        nent_o    => MPROJ_L3L4CD_L5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L5PHIC_AV_dout_mask
      );

    MPROJ_L3L4CD_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L5PHIC_wea,
        addra     => MPROJ_L3L4CD_L5PHIC_writeaddr,
        dina      => MPROJ_L3L4CD_L5PHIC_din,
        wea_out       => MPROJ_L3L4CD_L5PHIC_wea_delay,
        addra_out     => MPROJ_L3L4CD_L5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L5PHIC_start
      );

    MPROJ_L1L2G_L5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L5PHID_wea_delay,
        addra     => MPROJ_L1L2G_L5PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L5PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_L5PHID_V_dout,
        sync_nent => MPROJ_L1L2G_L5PHID_start,
        nent_o    => MPROJ_L1L2G_L5PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L5PHID_AV_dout_mask
      );

    MPROJ_L1L2G_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L5PHID_wea,
        addra     => MPROJ_L1L2G_L5PHID_writeaddr,
        dina      => MPROJ_L1L2G_L5PHID_din,
        wea_out       => MPROJ_L1L2G_L5PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_L5PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L5PHID_start
      );

    MPROJ_L1L2HI_L5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L5PHID_wea_delay,
        addra     => MPROJ_L1L2HI_L5PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L5PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_L5PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_L5PHID_start,
        nent_o    => MPROJ_L1L2HI_L5PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L5PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L5PHID_wea,
        addra     => MPROJ_L1L2HI_L5PHID_writeaddr,
        dina      => MPROJ_L1L2HI_L5PHID_din,
        wea_out       => MPROJ_L1L2HI_L5PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_L5PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L5PHID_start
      );

    MPROJ_L1L2JKL_L5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L5PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_L5PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L5PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L5PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_L5PHID_start,
        nent_o    => MPROJ_L1L2JKL_L5PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L5PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L5PHID_wea,
        addra     => MPROJ_L1L2JKL_L5PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_L5PHID_din,
        wea_out       => MPROJ_L1L2JKL_L5PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L5PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L5PHID_start
      );

    MPROJ_L2L3ABCD_L5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_L5PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_L5PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_L5PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_L5PHID_start,
        nent_o    => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_L5PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_L5PHID_wea,
        addra     => MPROJ_L2L3ABCD_L5PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_L5PHID_din,
        wea_out       => MPROJ_L2L3ABCD_L5PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_L5PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_L5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_L5PHID_start
      );

    MPROJ_L3L4CD_L5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L5PHID_wea_delay,
        addra     => MPROJ_L3L4CD_L5PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L5PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_L5PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_L5PHID_start,
        nent_o    => MPROJ_L3L4CD_L5PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L5PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L5PHID_wea,
        addra     => MPROJ_L3L4CD_L5PHID_writeaddr,
        dina      => MPROJ_L3L4CD_L5PHID_din,
        wea_out       => MPROJ_L3L4CD_L5PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_L5PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L5PHID_start
      );

    MPROJ_L1L2ABC_L6PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L6PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_L6PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L6PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L6PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_L6PHIA_start,
        nent_o    => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L6PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L6PHIA_wea,
        addra     => MPROJ_L1L2ABC_L6PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_L6PHIA_din,
        wea_out       => MPROJ_L1L2ABC_L6PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L6PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L6PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L6PHIA_start
      );

    MPROJ_L1L2DE_L6PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L6PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_L6PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L6PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_L6PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_L6PHIA_start,
        nent_o    => MPROJ_L1L2DE_L6PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L6PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L6PHIA_wea,
        addra     => MPROJ_L1L2DE_L6PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_L6PHIA_din,
        wea_out       => MPROJ_L1L2DE_L6PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_L6PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L6PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L6PHIA_start
      );

    MPROJ_L1L2F_L6PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L6PHIA_wea_delay,
        addra     => MPROJ_L1L2F_L6PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L6PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_L6PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_L6PHIA_start,
        nent_o    => MPROJ_L1L2F_L6PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L6PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L6PHIA_wea,
        addra     => MPROJ_L1L2F_L6PHIA_writeaddr,
        dina      => MPROJ_L1L2F_L6PHIA_din,
        wea_out       => MPROJ_L1L2F_L6PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_L6PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L6PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L6PHIA_start
      );

    MPROJ_L3L4AB_L6PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L6PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_L6PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L6PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_L6PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_L6PHIA_start,
        nent_o    => MPROJ_L3L4AB_L6PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L6PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L6PHIA_wea,
        addra     => MPROJ_L3L4AB_L6PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_L6PHIA_din,
        wea_out       => MPROJ_L3L4AB_L6PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_L6PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L6PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L6PHIA_start
      );

    MPROJ_L1L2ABC_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_L6PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_L6PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_L6PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_L6PHIB_start,
        nent_o    => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_L6PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_L6PHIB_wea,
        addra     => MPROJ_L1L2ABC_L6PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_L6PHIB_din,
        wea_out       => MPROJ_L1L2ABC_L6PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_L6PHIB_start
      );

    MPROJ_L1L2DE_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L6PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L6PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_L6PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_L6PHIB_start,
        nent_o    => MPROJ_L1L2DE_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L6PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L6PHIB_wea,
        addra     => MPROJ_L1L2DE_L6PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_L6PHIB_din,
        wea_out       => MPROJ_L1L2DE_L6PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L6PHIB_start
      );

    MPROJ_L1L2F_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L6PHIB_wea_delay,
        addra     => MPROJ_L1L2F_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L6PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_L6PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_L6PHIB_start,
        nent_o    => MPROJ_L1L2F_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L6PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L6PHIB_wea,
        addra     => MPROJ_L1L2F_L6PHIB_writeaddr,
        dina      => MPROJ_L1L2F_L6PHIB_din,
        wea_out       => MPROJ_L1L2F_L6PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L6PHIB_start
      );

    MPROJ_L1L2G_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L6PHIB_wea_delay,
        addra     => MPROJ_L1L2G_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L6PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_L6PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_L6PHIB_start,
        nent_o    => MPROJ_L1L2G_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L6PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L6PHIB_wea,
        addra     => MPROJ_L1L2G_L6PHIB_writeaddr,
        dina      => MPROJ_L1L2G_L6PHIB_din,
        wea_out       => MPROJ_L1L2G_L6PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L6PHIB_start
      );

    MPROJ_L1L2HI_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L6PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L6PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_L6PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_L6PHIB_start,
        nent_o    => MPROJ_L1L2HI_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L6PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L6PHIB_wea,
        addra     => MPROJ_L1L2HI_L6PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_L6PHIB_din,
        wea_out       => MPROJ_L1L2HI_L6PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L6PHIB_start
      );

    MPROJ_L3L4AB_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L6PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L6PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_L6PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_L6PHIB_start,
        nent_o    => MPROJ_L3L4AB_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L6PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L6PHIB_wea,
        addra     => MPROJ_L3L4AB_L6PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_L6PHIB_din,
        wea_out       => MPROJ_L3L4AB_L6PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L6PHIB_start
      );

    MPROJ_L3L4CD_L6PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L6PHIB_wea_delay,
        addra     => MPROJ_L3L4CD_L6PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L6PHIB_V_readaddr,
        doutb     => MPROJ_L3L4CD_L6PHIB_V_dout,
        sync_nent => MPROJ_L3L4CD_L6PHIB_start,
        nent_o    => MPROJ_L3L4CD_L6PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L6PHIB_AV_dout_mask
      );

    MPROJ_L3L4CD_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L6PHIB_wea,
        addra     => MPROJ_L3L4CD_L6PHIB_writeaddr,
        dina      => MPROJ_L3L4CD_L6PHIB_din,
        wea_out       => MPROJ_L3L4CD_L6PHIB_wea_delay,
        addra_out     => MPROJ_L3L4CD_L6PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L6PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L6PHIB_start
      );

    MPROJ_L1L2DE_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_L6PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_L6PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_L6PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_L6PHIC_start,
        nent_o    => MPROJ_L1L2DE_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_L6PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_L6PHIC_wea,
        addra     => MPROJ_L1L2DE_L6PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_L6PHIC_din,
        wea_out       => MPROJ_L1L2DE_L6PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_L6PHIC_start
      );

    MPROJ_L1L2F_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_L6PHIC_wea_delay,
        addra     => MPROJ_L1L2F_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_L6PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_L6PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_L6PHIC_start,
        nent_o    => MPROJ_L1L2F_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_L6PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_L6PHIC_wea,
        addra     => MPROJ_L1L2F_L6PHIC_writeaddr,
        dina      => MPROJ_L1L2F_L6PHIC_din,
        wea_out       => MPROJ_L1L2F_L6PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_L6PHIC_start
      );

    MPROJ_L1L2G_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L6PHIC_wea_delay,
        addra     => MPROJ_L1L2G_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L6PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_L6PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_L6PHIC_start,
        nent_o    => MPROJ_L1L2G_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L6PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L6PHIC_wea,
        addra     => MPROJ_L1L2G_L6PHIC_writeaddr,
        dina      => MPROJ_L1L2G_L6PHIC_din,
        wea_out       => MPROJ_L1L2G_L6PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L6PHIC_start
      );

    MPROJ_L1L2HI_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L6PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L6PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_L6PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_L6PHIC_start,
        nent_o    => MPROJ_L1L2HI_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L6PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L6PHIC_wea,
        addra     => MPROJ_L1L2HI_L6PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_L6PHIC_din,
        wea_out       => MPROJ_L1L2HI_L6PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L6PHIC_start
      );

    MPROJ_L1L2JKL_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L6PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L6PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L6PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_L6PHIC_start,
        nent_o    => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L6PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L6PHIC_wea,
        addra     => MPROJ_L1L2JKL_L6PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_L6PHIC_din,
        wea_out       => MPROJ_L1L2JKL_L6PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L6PHIC_start
      );

    MPROJ_L3L4AB_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_L6PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_L6PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_L6PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_L6PHIC_start,
        nent_o    => MPROJ_L3L4AB_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_L6PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_L6PHIC_wea,
        addra     => MPROJ_L3L4AB_L6PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_L6PHIC_din,
        wea_out       => MPROJ_L3L4AB_L6PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_L6PHIC_start
      );

    MPROJ_L3L4CD_L6PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L6PHIC_wea_delay,
        addra     => MPROJ_L3L4CD_L6PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L6PHIC_V_readaddr,
        doutb     => MPROJ_L3L4CD_L6PHIC_V_dout,
        sync_nent => MPROJ_L3L4CD_L6PHIC_start,
        nent_o    => MPROJ_L3L4CD_L6PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L6PHIC_AV_dout_mask
      );

    MPROJ_L3L4CD_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L6PHIC_wea,
        addra     => MPROJ_L3L4CD_L6PHIC_writeaddr,
        dina      => MPROJ_L3L4CD_L6PHIC_din,
        wea_out       => MPROJ_L3L4CD_L6PHIC_wea_delay,
        addra_out     => MPROJ_L3L4CD_L6PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L6PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L6PHIC_start
      );

    MPROJ_L1L2G_L6PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_L6PHID_wea_delay,
        addra     => MPROJ_L1L2G_L6PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_L6PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_L6PHID_V_dout,
        sync_nent => MPROJ_L1L2G_L6PHID_start,
        nent_o    => MPROJ_L1L2G_L6PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_L6PHID_AV_dout_mask
      );

    MPROJ_L1L2G_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_L6PHID_wea,
        addra     => MPROJ_L1L2G_L6PHID_writeaddr,
        dina      => MPROJ_L1L2G_L6PHID_din,
        wea_out       => MPROJ_L1L2G_L6PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_L6PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_L6PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_L6PHID_start
      );

    MPROJ_L1L2HI_L6PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_L6PHID_wea_delay,
        addra     => MPROJ_L1L2HI_L6PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_L6PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_L6PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_L6PHID_start,
        nent_o    => MPROJ_L1L2HI_L6PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_L6PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_L6PHID_wea,
        addra     => MPROJ_L1L2HI_L6PHID_writeaddr,
        dina      => MPROJ_L1L2HI_L6PHID_din,
        wea_out       => MPROJ_L1L2HI_L6PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_L6PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_L6PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_L6PHID_start
      );

    MPROJ_L1L2JKL_L6PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_L6PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_L6PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_L6PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_L6PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_L6PHID_start,
        nent_o    => MPROJ_L1L2JKL_L6PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_L6PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_L6PHID_wea,
        addra     => MPROJ_L1L2JKL_L6PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_L6PHID_din,
        wea_out       => MPROJ_L1L2JKL_L6PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_L6PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_L6PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_L6PHID_start
      );

    MPROJ_L3L4CD_L6PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_L6PHID_wea_delay,
        addra     => MPROJ_L3L4CD_L6PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_L6PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_L6PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_L6PHID_start,
        nent_o    => MPROJ_L3L4CD_L6PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_L6PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 58
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_L6PHID_wea,
        addra     => MPROJ_L3L4CD_L6PHID_writeaddr,
        dina      => MPROJ_L3L4CD_L6PHID_din,
        wea_out       => MPROJ_L3L4CD_L6PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_L6PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_L6PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_L6PHID_start
      );

    MPROJ_L1L2ABC_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D1PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_D1PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D1PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D1PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_D1PHIA_start,
        nent_o    => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D1PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D1PHIA_wea,
        addra     => MPROJ_L1L2ABC_D1PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_D1PHIA_din,
        wea_out       => MPROJ_L1L2ABC_D1PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D1PHIA_start
      );

    MPROJ_L1L2DE_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D1PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_D1PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D1PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_D1PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_D1PHIA_start,
        nent_o    => MPROJ_L1L2DE_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D1PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D1PHIA_wea,
        addra     => MPROJ_L1L2DE_D1PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_D1PHIA_din,
        wea_out       => MPROJ_L1L2DE_D1PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D1PHIA_start
      );

    MPROJ_L1L2F_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D1PHIA_wea_delay,
        addra     => MPROJ_L1L2F_D1PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D1PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_D1PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_D1PHIA_start,
        nent_o    => MPROJ_L1L2F_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D1PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D1PHIA_wea,
        addra     => MPROJ_L1L2F_D1PHIA_writeaddr,
        dina      => MPROJ_L1L2F_D1PHIA_din,
        wea_out       => MPROJ_L1L2F_D1PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D1PHIA_start
      );

    MPROJ_L2L3ABCD_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_D1PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D1PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D1PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D1PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D1PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIA_wea,
        addra     => MPROJ_L2L3ABCD_D1PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_D1PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_D1PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D1PHIA_start
      );

    MPROJ_L3L4AB_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D1PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_D1PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D1PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_D1PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_D1PHIA_start,
        nent_o    => MPROJ_L3L4AB_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D1PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D1PHIA_wea,
        addra     => MPROJ_L3L4AB_D1PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_D1PHIA_din,
        wea_out       => MPROJ_L3L4AB_D1PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D1PHIA_start
      );

    MPROJ_D3D4ABCD_D1PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIA_wea_delay,
        addra     => MPROJ_D3D4ABCD_D1PHIA_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D1PHIA_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D1PHIA_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D1PHIA_start,
        nent_o    => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D1PHIA_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIA_wea,
        addra     => MPROJ_D3D4ABCD_D1PHIA_writeaddr,
        dina      => MPROJ_D3D4ABCD_D1PHIA_din,
        wea_out       => MPROJ_D3D4ABCD_D1PHIA_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D1PHIA_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D1PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D1PHIA_start
      );

    MPROJ_L1L2ABC_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D1PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D1PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D1PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_D1PHIB_start,
        nent_o    => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D1PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D1PHIB_wea,
        addra     => MPROJ_L1L2ABC_D1PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_D1PHIB_din,
        wea_out       => MPROJ_L1L2ABC_D1PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D1PHIB_start
      );

    MPROJ_L1L2DE_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D1PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D1PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_D1PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_D1PHIB_start,
        nent_o    => MPROJ_L1L2DE_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D1PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D1PHIB_wea,
        addra     => MPROJ_L1L2DE_D1PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_D1PHIB_din,
        wea_out       => MPROJ_L1L2DE_D1PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D1PHIB_start
      );

    MPROJ_L1L2F_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D1PHIB_wea_delay,
        addra     => MPROJ_L1L2F_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D1PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_D1PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_D1PHIB_start,
        nent_o    => MPROJ_L1L2F_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D1PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D1PHIB_wea,
        addra     => MPROJ_L1L2F_D1PHIB_writeaddr,
        dina      => MPROJ_L1L2F_D1PHIB_din,
        wea_out       => MPROJ_L1L2F_D1PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D1PHIB_start
      );

    MPROJ_L1L2G_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D1PHIB_wea_delay,
        addra     => MPROJ_L1L2G_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D1PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_D1PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_D1PHIB_start,
        nent_o    => MPROJ_L1L2G_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D1PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D1PHIB_wea,
        addra     => MPROJ_L1L2G_D1PHIB_writeaddr,
        dina      => MPROJ_L1L2G_D1PHIB_din,
        wea_out       => MPROJ_L1L2G_D1PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D1PHIB_start
      );

    MPROJ_L1L2HI_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D1PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D1PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_D1PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_D1PHIB_start,
        nent_o    => MPROJ_L1L2HI_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D1PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D1PHIB_wea,
        addra     => MPROJ_L1L2HI_D1PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_D1PHIB_din,
        wea_out       => MPROJ_L1L2HI_D1PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D1PHIB_start
      );

    MPROJ_L2L3ABCD_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D1PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D1PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D1PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D1PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIB_wea,
        addra     => MPROJ_L2L3ABCD_D1PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_D1PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_D1PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D1PHIB_start
      );

    MPROJ_L3L4AB_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D1PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D1PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_D1PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_D1PHIB_start,
        nent_o    => MPROJ_L3L4AB_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D1PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D1PHIB_wea,
        addra     => MPROJ_L3L4AB_D1PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_D1PHIB_din,
        wea_out       => MPROJ_L3L4AB_D1PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D1PHIB_start
      );

    MPROJ_L3L4CD_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D1PHIB_wea_delay,
        addra     => MPROJ_L3L4CD_D1PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D1PHIB_V_readaddr,
        doutb     => MPROJ_L3L4CD_D1PHIB_V_dout,
        sync_nent => MPROJ_L3L4CD_D1PHIB_start,
        nent_o    => MPROJ_L3L4CD_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D1PHIB_AV_dout_mask
      );

    MPROJ_L3L4CD_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D1PHIB_wea,
        addra     => MPROJ_L3L4CD_D1PHIB_writeaddr,
        dina      => MPROJ_L3L4CD_D1PHIB_din,
        wea_out       => MPROJ_L3L4CD_D1PHIB_wea_delay,
        addra_out     => MPROJ_L3L4CD_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D1PHIB_start
      );

    MPROJ_D3D4ABCD_D1PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIB_wea_delay,
        addra     => MPROJ_D3D4ABCD_D1PHIB_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D1PHIB_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D1PHIB_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D1PHIB_start,
        nent_o    => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D1PHIB_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIB_wea,
        addra     => MPROJ_D3D4ABCD_D1PHIB_writeaddr,
        dina      => MPROJ_D3D4ABCD_D1PHIB_din,
        wea_out       => MPROJ_D3D4ABCD_D1PHIB_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D1PHIB_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D1PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D1PHIB_start
      );

    MPROJ_L1L2DE_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D1PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D1PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_D1PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_D1PHIC_start,
        nent_o    => MPROJ_L1L2DE_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D1PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D1PHIC_wea,
        addra     => MPROJ_L1L2DE_D1PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_D1PHIC_din,
        wea_out       => MPROJ_L1L2DE_D1PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D1PHIC_start
      );

    MPROJ_L1L2F_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D1PHIC_wea_delay,
        addra     => MPROJ_L1L2F_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D1PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_D1PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_D1PHIC_start,
        nent_o    => MPROJ_L1L2F_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D1PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D1PHIC_wea,
        addra     => MPROJ_L1L2F_D1PHIC_writeaddr,
        dina      => MPROJ_L1L2F_D1PHIC_din,
        wea_out       => MPROJ_L1L2F_D1PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D1PHIC_start
      );

    MPROJ_L1L2G_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D1PHIC_wea_delay,
        addra     => MPROJ_L1L2G_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D1PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_D1PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_D1PHIC_start,
        nent_o    => MPROJ_L1L2G_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D1PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D1PHIC_wea,
        addra     => MPROJ_L1L2G_D1PHIC_writeaddr,
        dina      => MPROJ_L1L2G_D1PHIC_din,
        wea_out       => MPROJ_L1L2G_D1PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D1PHIC_start
      );

    MPROJ_L1L2HI_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D1PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D1PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_D1PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_D1PHIC_start,
        nent_o    => MPROJ_L1L2HI_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D1PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D1PHIC_wea,
        addra     => MPROJ_L1L2HI_D1PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_D1PHIC_din,
        wea_out       => MPROJ_L1L2HI_D1PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D1PHIC_start
      );

    MPROJ_L1L2JKL_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D1PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D1PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D1PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_D1PHIC_start,
        nent_o    => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D1PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D1PHIC_wea,
        addra     => MPROJ_L1L2JKL_D1PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_D1PHIC_din,
        wea_out       => MPROJ_L1L2JKL_D1PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D1PHIC_start
      );

    MPROJ_L2L3ABCD_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D1PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D1PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D1PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D1PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHIC_wea,
        addra     => MPROJ_L2L3ABCD_D1PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_D1PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_D1PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D1PHIC_start
      );

    MPROJ_L3L4AB_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D1PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D1PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_D1PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_D1PHIC_start,
        nent_o    => MPROJ_L3L4AB_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D1PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D1PHIC_wea,
        addra     => MPROJ_L3L4AB_D1PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_D1PHIC_din,
        wea_out       => MPROJ_L3L4AB_D1PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D1PHIC_start
      );

    MPROJ_L3L4CD_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D1PHIC_wea_delay,
        addra     => MPROJ_L3L4CD_D1PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D1PHIC_V_readaddr,
        doutb     => MPROJ_L3L4CD_D1PHIC_V_dout,
        sync_nent => MPROJ_L3L4CD_D1PHIC_start,
        nent_o    => MPROJ_L3L4CD_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D1PHIC_AV_dout_mask
      );

    MPROJ_L3L4CD_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D1PHIC_wea,
        addra     => MPROJ_L3L4CD_D1PHIC_writeaddr,
        dina      => MPROJ_L3L4CD_D1PHIC_din,
        wea_out       => MPROJ_L3L4CD_D1PHIC_wea_delay,
        addra_out     => MPROJ_L3L4CD_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D1PHIC_start
      );

    MPROJ_D3D4ABCD_D1PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIC_wea_delay,
        addra     => MPROJ_D3D4ABCD_D1PHIC_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D1PHIC_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D1PHIC_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D1PHIC_start,
        nent_o    => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D1PHIC_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHIC_wea,
        addra     => MPROJ_D3D4ABCD_D1PHIC_writeaddr,
        dina      => MPROJ_D3D4ABCD_D1PHIC_din,
        wea_out       => MPROJ_D3D4ABCD_D1PHIC_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D1PHIC_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D1PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D1PHIC_start
      );

    MPROJ_L1L2G_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D1PHID_wea_delay,
        addra     => MPROJ_L1L2G_D1PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D1PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_D1PHID_V_dout,
        sync_nent => MPROJ_L1L2G_D1PHID_start,
        nent_o    => MPROJ_L1L2G_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D1PHID_AV_dout_mask
      );

    MPROJ_L1L2G_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D1PHID_wea,
        addra     => MPROJ_L1L2G_D1PHID_writeaddr,
        dina      => MPROJ_L1L2G_D1PHID_din,
        wea_out       => MPROJ_L1L2G_D1PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D1PHID_start
      );

    MPROJ_L1L2HI_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D1PHID_wea_delay,
        addra     => MPROJ_L1L2HI_D1PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D1PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_D1PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_D1PHID_start,
        nent_o    => MPROJ_L1L2HI_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D1PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D1PHID_wea,
        addra     => MPROJ_L1L2HI_D1PHID_writeaddr,
        dina      => MPROJ_L1L2HI_D1PHID_din,
        wea_out       => MPROJ_L1L2HI_D1PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D1PHID_start
      );

    MPROJ_L1L2JKL_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D1PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_D1PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D1PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D1PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_D1PHID_start,
        nent_o    => MPROJ_L1L2JKL_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D1PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D1PHID_wea,
        addra     => MPROJ_L1L2JKL_D1PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_D1PHID_din,
        wea_out       => MPROJ_L1L2JKL_D1PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D1PHID_start
      );

    MPROJ_L2L3ABCD_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_D1PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D1PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D1PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D1PHID_start,
        nent_o    => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D1PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D1PHID_wea,
        addra     => MPROJ_L2L3ABCD_D1PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_D1PHID_din,
        wea_out       => MPROJ_L2L3ABCD_D1PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D1PHID_start
      );

    MPROJ_L3L4CD_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D1PHID_wea_delay,
        addra     => MPROJ_L3L4CD_D1PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D1PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_D1PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_D1PHID_start,
        nent_o    => MPROJ_L3L4CD_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D1PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D1PHID_wea,
        addra     => MPROJ_L3L4CD_D1PHID_writeaddr,
        dina      => MPROJ_L3L4CD_D1PHID_din,
        wea_out       => MPROJ_L3L4CD_D1PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D1PHID_start
      );

    MPROJ_D3D4ABCD_D1PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHID_wea_delay,
        addra     => MPROJ_D3D4ABCD_D1PHID_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D1PHID_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D1PHID_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D1PHID_start,
        nent_o    => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D1PHID_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D1PHID_wea,
        addra     => MPROJ_D3D4ABCD_D1PHID_writeaddr,
        dina      => MPROJ_D3D4ABCD_D1PHID_din,
        wea_out       => MPROJ_D3D4ABCD_D1PHID_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D1PHID_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D1PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D1PHID_start
      );

    MPROJ_L1L2ABC_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D2PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D2PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D2PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_D2PHIA_start,
        nent_o    => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D2PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D2PHIA_wea,
        addra     => MPROJ_L1L2ABC_D2PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_D2PHIA_din,
        wea_out       => MPROJ_L1L2ABC_D2PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D2PHIA_start
      );

    MPROJ_L1L2DE_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D2PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D2PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_D2PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_D2PHIA_start,
        nent_o    => MPROJ_L1L2DE_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D2PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D2PHIA_wea,
        addra     => MPROJ_L1L2DE_D2PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_D2PHIA_din,
        wea_out       => MPROJ_L1L2DE_D2PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D2PHIA_start
      );

    MPROJ_L1L2F_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D2PHIA_wea_delay,
        addra     => MPROJ_L1L2F_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D2PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_D2PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_D2PHIA_start,
        nent_o    => MPROJ_L1L2F_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D2PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D2PHIA_wea,
        addra     => MPROJ_L1L2F_D2PHIA_writeaddr,
        dina      => MPROJ_L1L2F_D2PHIA_din,
        wea_out       => MPROJ_L1L2F_D2PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D2PHIA_start
      );

    MPROJ_L2L3ABCD_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D2PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D2PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D2PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D2PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIA_wea,
        addra     => MPROJ_L2L3ABCD_D2PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_D2PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_D2PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D2PHIA_start
      );

    MPROJ_L3L4AB_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D2PHIA_wea_delay,
        addra     => MPROJ_L3L4AB_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D2PHIA_V_readaddr,
        doutb     => MPROJ_L3L4AB_D2PHIA_V_dout,
        sync_nent => MPROJ_L3L4AB_D2PHIA_start,
        nent_o    => MPROJ_L3L4AB_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D2PHIA_AV_dout_mask
      );

    MPROJ_L3L4AB_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D2PHIA_wea,
        addra     => MPROJ_L3L4AB_D2PHIA_writeaddr,
        dina      => MPROJ_L3L4AB_D2PHIA_din,
        wea_out       => MPROJ_L3L4AB_D2PHIA_wea_delay,
        addra_out     => MPROJ_L3L4AB_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D2PHIA_start
      );

    MPROJ_D3D4ABCD_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIA_wea_delay,
        addra     => MPROJ_D3D4ABCD_D2PHIA_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D2PHIA_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D2PHIA_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D2PHIA_start,
        nent_o    => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D2PHIA_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIA_wea,
        addra     => MPROJ_D3D4ABCD_D2PHIA_writeaddr,
        dina      => MPROJ_D3D4ABCD_D2PHIA_din,
        wea_out       => MPROJ_D3D4ABCD_D2PHIA_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D2PHIA_start
      );

    MPROJ_L1D1ABCD_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIA_wea_delay,
        addra     => MPROJ_L1D1ABCD_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D2PHIA_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D2PHIA_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D2PHIA_start,
        nent_o    => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D2PHIA_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIA_wea,
        addra     => MPROJ_L1D1ABCD_D2PHIA_writeaddr,
        dina      => MPROJ_L1D1ABCD_D2PHIA_din,
        wea_out       => MPROJ_L1D1ABCD_D2PHIA_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D2PHIA_start
      );

    MPROJ_L2D1ABCD_D2PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIA_wea_delay,
        addra     => MPROJ_L2D1ABCD_D2PHIA_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D2PHIA_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D2PHIA_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D2PHIA_start,
        nent_o    => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D2PHIA_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIA_wea,
        addra     => MPROJ_L2D1ABCD_D2PHIA_writeaddr,
        dina      => MPROJ_L2D1ABCD_D2PHIA_din,
        wea_out       => MPROJ_L2D1ABCD_D2PHIA_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D2PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D2PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D2PHIA_start
      );

    MPROJ_L1L2ABC_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D2PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D2PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_D2PHIB_start,
        nent_o    => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D2PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D2PHIB_wea,
        addra     => MPROJ_L1L2ABC_D2PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_D2PHIB_din,
        wea_out       => MPROJ_L1L2ABC_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D2PHIB_start
      );

    MPROJ_L1L2DE_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D2PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_D2PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_D2PHIB_start,
        nent_o    => MPROJ_L1L2DE_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D2PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D2PHIB_wea,
        addra     => MPROJ_L1L2DE_D2PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_D2PHIB_din,
        wea_out       => MPROJ_L1L2DE_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D2PHIB_start
      );

    MPROJ_L1L2F_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D2PHIB_wea_delay,
        addra     => MPROJ_L1L2F_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_D2PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_D2PHIB_start,
        nent_o    => MPROJ_L1L2F_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D2PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D2PHIB_wea,
        addra     => MPROJ_L1L2F_D2PHIB_writeaddr,
        dina      => MPROJ_L1L2F_D2PHIB_din,
        wea_out       => MPROJ_L1L2F_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D2PHIB_start
      );

    MPROJ_L1L2G_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D2PHIB_wea_delay,
        addra     => MPROJ_L1L2G_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_D2PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_D2PHIB_start,
        nent_o    => MPROJ_L1L2G_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D2PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D2PHIB_wea,
        addra     => MPROJ_L1L2G_D2PHIB_writeaddr,
        dina      => MPROJ_L1L2G_D2PHIB_din,
        wea_out       => MPROJ_L1L2G_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D2PHIB_start
      );

    MPROJ_L1L2HI_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D2PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_D2PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_D2PHIB_start,
        nent_o    => MPROJ_L1L2HI_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D2PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D2PHIB_wea,
        addra     => MPROJ_L1L2HI_D2PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_D2PHIB_din,
        wea_out       => MPROJ_L1L2HI_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D2PHIB_start
      );

    MPROJ_L2L3ABCD_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D2PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D2PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D2PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D2PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIB_wea,
        addra     => MPROJ_L2L3ABCD_D2PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_D2PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_D2PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D2PHIB_start
      );

    MPROJ_L3L4AB_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D2PHIB_wea_delay,
        addra     => MPROJ_L3L4AB_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D2PHIB_V_readaddr,
        doutb     => MPROJ_L3L4AB_D2PHIB_V_dout,
        sync_nent => MPROJ_L3L4AB_D2PHIB_start,
        nent_o    => MPROJ_L3L4AB_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D2PHIB_AV_dout_mask
      );

    MPROJ_L3L4AB_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D2PHIB_wea,
        addra     => MPROJ_L3L4AB_D2PHIB_writeaddr,
        dina      => MPROJ_L3L4AB_D2PHIB_din,
        wea_out       => MPROJ_L3L4AB_D2PHIB_wea_delay,
        addra_out     => MPROJ_L3L4AB_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D2PHIB_start
      );

    MPROJ_L3L4CD_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D2PHIB_wea_delay,
        addra     => MPROJ_L3L4CD_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D2PHIB_V_readaddr,
        doutb     => MPROJ_L3L4CD_D2PHIB_V_dout,
        sync_nent => MPROJ_L3L4CD_D2PHIB_start,
        nent_o    => MPROJ_L3L4CD_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D2PHIB_AV_dout_mask
      );

    MPROJ_L3L4CD_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D2PHIB_wea,
        addra     => MPROJ_L3L4CD_D2PHIB_writeaddr,
        dina      => MPROJ_L3L4CD_D2PHIB_din,
        wea_out       => MPROJ_L3L4CD_D2PHIB_wea_delay,
        addra_out     => MPROJ_L3L4CD_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D2PHIB_start
      );

    MPROJ_D3D4ABCD_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIB_wea_delay,
        addra     => MPROJ_D3D4ABCD_D2PHIB_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D2PHIB_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D2PHIB_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D2PHIB_start,
        nent_o    => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D2PHIB_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIB_wea,
        addra     => MPROJ_D3D4ABCD_D2PHIB_writeaddr,
        dina      => MPROJ_D3D4ABCD_D2PHIB_din,
        wea_out       => MPROJ_D3D4ABCD_D2PHIB_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D2PHIB_start
      );

    MPROJ_L1D1ABCD_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIB_wea_delay,
        addra     => MPROJ_L1D1ABCD_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D2PHIB_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D2PHIB_start,
        nent_o    => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D2PHIB_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIB_wea,
        addra     => MPROJ_L1D1ABCD_D2PHIB_writeaddr,
        dina      => MPROJ_L1D1ABCD_D2PHIB_din,
        wea_out       => MPROJ_L1D1ABCD_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D2PHIB_start
      );

    MPROJ_L1D1EFGH_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHIB_wea_delay,
        addra     => MPROJ_L1D1EFGH_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D2PHIB_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D2PHIB_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D2PHIB_start,
        nent_o    => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D2PHIB_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHIB_wea,
        addra     => MPROJ_L1D1EFGH_D2PHIB_writeaddr,
        dina      => MPROJ_L1D1EFGH_D2PHIB_din,
        wea_out       => MPROJ_L1D1EFGH_D2PHIB_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D2PHIB_start
      );

    MPROJ_L2D1ABCD_D2PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIB_wea_delay,
        addra     => MPROJ_L2D1ABCD_D2PHIB_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D2PHIB_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D2PHIB_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D2PHIB_start,
        nent_o    => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D2PHIB_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIB_wea,
        addra     => MPROJ_L2D1ABCD_D2PHIB_writeaddr,
        dina      => MPROJ_L2D1ABCD_D2PHIB_din,
        wea_out       => MPROJ_L2D1ABCD_D2PHIB_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D2PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D2PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D2PHIB_start
      );

    MPROJ_L1L2DE_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D2PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_D2PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_D2PHIC_start,
        nent_o    => MPROJ_L1L2DE_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D2PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D2PHIC_wea,
        addra     => MPROJ_L1L2DE_D2PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_D2PHIC_din,
        wea_out       => MPROJ_L1L2DE_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D2PHIC_start
      );

    MPROJ_L1L2F_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D2PHIC_wea_delay,
        addra     => MPROJ_L1L2F_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_D2PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_D2PHIC_start,
        nent_o    => MPROJ_L1L2F_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D2PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D2PHIC_wea,
        addra     => MPROJ_L1L2F_D2PHIC_writeaddr,
        dina      => MPROJ_L1L2F_D2PHIC_din,
        wea_out       => MPROJ_L1L2F_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D2PHIC_start
      );

    MPROJ_L1L2G_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D2PHIC_wea_delay,
        addra     => MPROJ_L1L2G_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_D2PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_D2PHIC_start,
        nent_o    => MPROJ_L1L2G_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D2PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D2PHIC_wea,
        addra     => MPROJ_L1L2G_D2PHIC_writeaddr,
        dina      => MPROJ_L1L2G_D2PHIC_din,
        wea_out       => MPROJ_L1L2G_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D2PHIC_start
      );

    MPROJ_L1L2HI_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D2PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_D2PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_D2PHIC_start,
        nent_o    => MPROJ_L1L2HI_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D2PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D2PHIC_wea,
        addra     => MPROJ_L1L2HI_D2PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_D2PHIC_din,
        wea_out       => MPROJ_L1L2HI_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D2PHIC_start
      );

    MPROJ_L1L2JKL_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D2PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D2PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_D2PHIC_start,
        nent_o    => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D2PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D2PHIC_wea,
        addra     => MPROJ_L1L2JKL_D2PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_D2PHIC_din,
        wea_out       => MPROJ_L1L2JKL_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D2PHIC_start
      );

    MPROJ_L2L3ABCD_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D2PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D2PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D2PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D2PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHIC_wea,
        addra     => MPROJ_L2L3ABCD_D2PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_D2PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_D2PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D2PHIC_start
      );

    MPROJ_L3L4AB_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4AB_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4AB_D2PHIC_wea_delay,
        addra     => MPROJ_L3L4AB_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4AB_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4AB_D2PHIC_V_readaddr,
        doutb     => MPROJ_L3L4AB_D2PHIC_V_dout,
        sync_nent => MPROJ_L3L4AB_D2PHIC_start,
        nent_o    => MPROJ_L3L4AB_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4AB_D2PHIC_AV_dout_mask
      );

    MPROJ_L3L4AB_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4AB_D2PHIC_wea,
        addra     => MPROJ_L3L4AB_D2PHIC_writeaddr,
        dina      => MPROJ_L3L4AB_D2PHIC_din,
        wea_out       => MPROJ_L3L4AB_D2PHIC_wea_delay,
        addra_out     => MPROJ_L3L4AB_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4AB_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4AB_D2PHIC_start
      );

    MPROJ_L3L4CD_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D2PHIC_wea_delay,
        addra     => MPROJ_L3L4CD_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D2PHIC_V_readaddr,
        doutb     => MPROJ_L3L4CD_D2PHIC_V_dout,
        sync_nent => MPROJ_L3L4CD_D2PHIC_start,
        nent_o    => MPROJ_L3L4CD_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D2PHIC_AV_dout_mask
      );

    MPROJ_L3L4CD_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D2PHIC_wea,
        addra     => MPROJ_L3L4CD_D2PHIC_writeaddr,
        dina      => MPROJ_L3L4CD_D2PHIC_din,
        wea_out       => MPROJ_L3L4CD_D2PHIC_wea_delay,
        addra_out     => MPROJ_L3L4CD_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D2PHIC_start
      );

    MPROJ_D3D4ABCD_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIC_wea_delay,
        addra     => MPROJ_D3D4ABCD_D2PHIC_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D2PHIC_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D2PHIC_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D2PHIC_start,
        nent_o    => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D2PHIC_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHIC_wea,
        addra     => MPROJ_D3D4ABCD_D2PHIC_writeaddr,
        dina      => MPROJ_D3D4ABCD_D2PHIC_din,
        wea_out       => MPROJ_D3D4ABCD_D2PHIC_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D2PHIC_start
      );

    MPROJ_L1D1ABCD_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIC_wea_delay,
        addra     => MPROJ_L1D1ABCD_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D2PHIC_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D2PHIC_start,
        nent_o    => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D2PHIC_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D2PHIC_wea,
        addra     => MPROJ_L1D1ABCD_D2PHIC_writeaddr,
        dina      => MPROJ_L1D1ABCD_D2PHIC_din,
        wea_out       => MPROJ_L1D1ABCD_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D2PHIC_start
      );

    MPROJ_L1D1EFGH_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHIC_wea_delay,
        addra     => MPROJ_L1D1EFGH_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D2PHIC_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D2PHIC_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D2PHIC_start,
        nent_o    => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D2PHIC_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHIC_wea,
        addra     => MPROJ_L1D1EFGH_D2PHIC_writeaddr,
        dina      => MPROJ_L1D1EFGH_D2PHIC_din,
        wea_out       => MPROJ_L1D1EFGH_D2PHIC_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D2PHIC_start
      );

    MPROJ_L2D1ABCD_D2PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIC_wea_delay,
        addra     => MPROJ_L2D1ABCD_D2PHIC_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D2PHIC_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D2PHIC_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D2PHIC_start,
        nent_o    => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D2PHIC_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHIC_wea,
        addra     => MPROJ_L2D1ABCD_D2PHIC_writeaddr,
        dina      => MPROJ_L2D1ABCD_D2PHIC_din,
        wea_out       => MPROJ_L2D1ABCD_D2PHIC_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D2PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D2PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D2PHIC_start
      );

    MPROJ_L1L2G_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D2PHID_wea_delay,
        addra     => MPROJ_L1L2G_D2PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D2PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_D2PHID_V_dout,
        sync_nent => MPROJ_L1L2G_D2PHID_start,
        nent_o    => MPROJ_L1L2G_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D2PHID_AV_dout_mask
      );

    MPROJ_L1L2G_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D2PHID_wea,
        addra     => MPROJ_L1L2G_D2PHID_writeaddr,
        dina      => MPROJ_L1L2G_D2PHID_din,
        wea_out       => MPROJ_L1L2G_D2PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D2PHID_start
      );

    MPROJ_L1L2HI_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D2PHID_wea_delay,
        addra     => MPROJ_L1L2HI_D2PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D2PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_D2PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_D2PHID_start,
        nent_o    => MPROJ_L1L2HI_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D2PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D2PHID_wea,
        addra     => MPROJ_L1L2HI_D2PHID_writeaddr,
        dina      => MPROJ_L1L2HI_D2PHID_din,
        wea_out       => MPROJ_L1L2HI_D2PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D2PHID_start
      );

    MPROJ_L1L2JKL_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D2PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_D2PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D2PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D2PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_D2PHID_start,
        nent_o    => MPROJ_L1L2JKL_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D2PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D2PHID_wea,
        addra     => MPROJ_L1L2JKL_D2PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_D2PHID_din,
        wea_out       => MPROJ_L1L2JKL_D2PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D2PHID_start
      );

    MPROJ_L2L3ABCD_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_D2PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D2PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D2PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D2PHID_start,
        nent_o    => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D2PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D2PHID_wea,
        addra     => MPROJ_L2L3ABCD_D2PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_D2PHID_din,
        wea_out       => MPROJ_L2L3ABCD_D2PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D2PHID_start
      );

    MPROJ_L3L4CD_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L3L4CD_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L3L4CD_D2PHID_wea_delay,
        addra     => MPROJ_L3L4CD_D2PHID_writeaddr_delay,
        dina      => MPROJ_L3L4CD_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L3L4CD_D2PHID_V_readaddr,
        doutb     => MPROJ_L3L4CD_D2PHID_V_dout,
        sync_nent => MPROJ_L3L4CD_D2PHID_start,
        nent_o    => MPROJ_L3L4CD_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L3L4CD_D2PHID_AV_dout_mask
      );

    MPROJ_L3L4CD_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L3L4CD_D2PHID_wea,
        addra     => MPROJ_L3L4CD_D2PHID_writeaddr,
        dina      => MPROJ_L3L4CD_D2PHID_din,
        wea_out       => MPROJ_L3L4CD_D2PHID_wea_delay,
        addra_out     => MPROJ_L3L4CD_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L3L4CD_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L3L4CD_D2PHID_start
      );

    MPROJ_D3D4ABCD_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHID_wea_delay,
        addra     => MPROJ_D3D4ABCD_D2PHID_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D2PHID_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D2PHID_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D2PHID_start,
        nent_o    => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D2PHID_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D2PHID_wea,
        addra     => MPROJ_D3D4ABCD_D2PHID_writeaddr,
        dina      => MPROJ_D3D4ABCD_D2PHID_din,
        wea_out       => MPROJ_D3D4ABCD_D2PHID_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D2PHID_start
      );

    MPROJ_L1D1EFGH_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHID_wea_delay,
        addra     => MPROJ_L1D1EFGH_D2PHID_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D2PHID_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D2PHID_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D2PHID_start,
        nent_o    => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D2PHID_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D2PHID_wea,
        addra     => MPROJ_L1D1EFGH_D2PHID_writeaddr,
        dina      => MPROJ_L1D1EFGH_D2PHID_din,
        wea_out       => MPROJ_L1D1EFGH_D2PHID_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D2PHID_start
      );

    MPROJ_L2D1ABCD_D2PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHID_wea_delay,
        addra     => MPROJ_L2D1ABCD_D2PHID_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D2PHID_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D2PHID_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D2PHID_start,
        nent_o    => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D2PHID_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D2PHID_wea,
        addra     => MPROJ_L2D1ABCD_D2PHID_writeaddr,
        dina      => MPROJ_L2D1ABCD_D2PHID_din,
        wea_out       => MPROJ_L2D1ABCD_D2PHID_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D2PHID_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D2PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D2PHID_start
      );

    MPROJ_L1L2ABC_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D3PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D3PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D3PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_D3PHIA_start,
        nent_o    => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D3PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D3PHIA_wea,
        addra     => MPROJ_L1L2ABC_D3PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_D3PHIA_din,
        wea_out       => MPROJ_L1L2ABC_D3PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D3PHIA_start
      );

    MPROJ_L1L2DE_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D3PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D3PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_D3PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_D3PHIA_start,
        nent_o    => MPROJ_L1L2DE_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D3PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D3PHIA_wea,
        addra     => MPROJ_L1L2DE_D3PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_D3PHIA_din,
        wea_out       => MPROJ_L1L2DE_D3PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D3PHIA_start
      );

    MPROJ_L1L2F_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D3PHIA_wea_delay,
        addra     => MPROJ_L1L2F_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D3PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_D3PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_D3PHIA_start,
        nent_o    => MPROJ_L1L2F_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D3PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D3PHIA_wea,
        addra     => MPROJ_L1L2F_D3PHIA_writeaddr,
        dina      => MPROJ_L1L2F_D3PHIA_din,
        wea_out       => MPROJ_L1L2F_D3PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D3PHIA_start
      );

    MPROJ_L2L3ABCD_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D3PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D3PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D3PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D3PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIA_wea,
        addra     => MPROJ_L2L3ABCD_D3PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_D3PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_D3PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D3PHIA_start
      );

    MPROJ_D1D2ABCD_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIA_wea_delay,
        addra     => MPROJ_D1D2ABCD_D3PHIA_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D3PHIA_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D3PHIA_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D3PHIA_start,
        nent_o    => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D3PHIA_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIA_wea,
        addra     => MPROJ_D1D2ABCD_D3PHIA_writeaddr,
        dina      => MPROJ_D1D2ABCD_D3PHIA_din,
        wea_out       => MPROJ_D1D2ABCD_D3PHIA_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D3PHIA_start
      );

    MPROJ_L1D1ABCD_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIA_wea_delay,
        addra     => MPROJ_L1D1ABCD_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D3PHIA_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D3PHIA_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D3PHIA_start,
        nent_o    => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D3PHIA_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIA_wea,
        addra     => MPROJ_L1D1ABCD_D3PHIA_writeaddr,
        dina      => MPROJ_L1D1ABCD_D3PHIA_din,
        wea_out       => MPROJ_L1D1ABCD_D3PHIA_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D3PHIA_start
      );

    MPROJ_L2D1ABCD_D3PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIA_wea_delay,
        addra     => MPROJ_L2D1ABCD_D3PHIA_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D3PHIA_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D3PHIA_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D3PHIA_start,
        nent_o    => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D3PHIA_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIA_wea,
        addra     => MPROJ_L2D1ABCD_D3PHIA_writeaddr,
        dina      => MPROJ_L2D1ABCD_D3PHIA_din,
        wea_out       => MPROJ_L2D1ABCD_D3PHIA_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D3PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D3PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D3PHIA_start
      );

    MPROJ_L1L2ABC_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D3PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D3PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_D3PHIB_start,
        nent_o    => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D3PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D3PHIB_wea,
        addra     => MPROJ_L1L2ABC_D3PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_D3PHIB_din,
        wea_out       => MPROJ_L1L2ABC_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D3PHIB_start
      );

    MPROJ_L1L2DE_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D3PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_D3PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_D3PHIB_start,
        nent_o    => MPROJ_L1L2DE_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D3PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D3PHIB_wea,
        addra     => MPROJ_L1L2DE_D3PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_D3PHIB_din,
        wea_out       => MPROJ_L1L2DE_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D3PHIB_start
      );

    MPROJ_L1L2F_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D3PHIB_wea_delay,
        addra     => MPROJ_L1L2F_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_D3PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_D3PHIB_start,
        nent_o    => MPROJ_L1L2F_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D3PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D3PHIB_wea,
        addra     => MPROJ_L1L2F_D3PHIB_writeaddr,
        dina      => MPROJ_L1L2F_D3PHIB_din,
        wea_out       => MPROJ_L1L2F_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D3PHIB_start
      );

    MPROJ_L1L2G_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D3PHIB_wea_delay,
        addra     => MPROJ_L1L2G_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_D3PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_D3PHIB_start,
        nent_o    => MPROJ_L1L2G_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D3PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D3PHIB_wea,
        addra     => MPROJ_L1L2G_D3PHIB_writeaddr,
        dina      => MPROJ_L1L2G_D3PHIB_din,
        wea_out       => MPROJ_L1L2G_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D3PHIB_start
      );

    MPROJ_L1L2HI_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D3PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_D3PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_D3PHIB_start,
        nent_o    => MPROJ_L1L2HI_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D3PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D3PHIB_wea,
        addra     => MPROJ_L1L2HI_D3PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_D3PHIB_din,
        wea_out       => MPROJ_L1L2HI_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D3PHIB_start
      );

    MPROJ_L2L3ABCD_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D3PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D3PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D3PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D3PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIB_wea,
        addra     => MPROJ_L2L3ABCD_D3PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_D3PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_D3PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D3PHIB_start
      );

    MPROJ_D1D2ABCD_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIB_wea_delay,
        addra     => MPROJ_D1D2ABCD_D3PHIB_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D3PHIB_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D3PHIB_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D3PHIB_start,
        nent_o    => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D3PHIB_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIB_wea,
        addra     => MPROJ_D1D2ABCD_D3PHIB_writeaddr,
        dina      => MPROJ_D1D2ABCD_D3PHIB_din,
        wea_out       => MPROJ_D1D2ABCD_D3PHIB_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D3PHIB_start
      );

    MPROJ_L1D1ABCD_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIB_wea_delay,
        addra     => MPROJ_L1D1ABCD_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D3PHIB_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D3PHIB_start,
        nent_o    => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D3PHIB_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIB_wea,
        addra     => MPROJ_L1D1ABCD_D3PHIB_writeaddr,
        dina      => MPROJ_L1D1ABCD_D3PHIB_din,
        wea_out       => MPROJ_L1D1ABCD_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D3PHIB_start
      );

    MPROJ_L1D1EFGH_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHIB_wea_delay,
        addra     => MPROJ_L1D1EFGH_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D3PHIB_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D3PHIB_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D3PHIB_start,
        nent_o    => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D3PHIB_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHIB_wea,
        addra     => MPROJ_L1D1EFGH_D3PHIB_writeaddr,
        dina      => MPROJ_L1D1EFGH_D3PHIB_din,
        wea_out       => MPROJ_L1D1EFGH_D3PHIB_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D3PHIB_start
      );

    MPROJ_L2D1ABCD_D3PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIB_wea_delay,
        addra     => MPROJ_L2D1ABCD_D3PHIB_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D3PHIB_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D3PHIB_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D3PHIB_start,
        nent_o    => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D3PHIB_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIB_wea,
        addra     => MPROJ_L2D1ABCD_D3PHIB_writeaddr,
        dina      => MPROJ_L2D1ABCD_D3PHIB_din,
        wea_out       => MPROJ_L2D1ABCD_D3PHIB_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D3PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D3PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D3PHIB_start
      );

    MPROJ_L1L2DE_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D3PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_D3PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_D3PHIC_start,
        nent_o    => MPROJ_L1L2DE_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D3PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D3PHIC_wea,
        addra     => MPROJ_L1L2DE_D3PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_D3PHIC_din,
        wea_out       => MPROJ_L1L2DE_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D3PHIC_start
      );

    MPROJ_L1L2F_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D3PHIC_wea_delay,
        addra     => MPROJ_L1L2F_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_D3PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_D3PHIC_start,
        nent_o    => MPROJ_L1L2F_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D3PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D3PHIC_wea,
        addra     => MPROJ_L1L2F_D3PHIC_writeaddr,
        dina      => MPROJ_L1L2F_D3PHIC_din,
        wea_out       => MPROJ_L1L2F_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D3PHIC_start
      );

    MPROJ_L1L2G_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D3PHIC_wea_delay,
        addra     => MPROJ_L1L2G_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_D3PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_D3PHIC_start,
        nent_o    => MPROJ_L1L2G_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D3PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D3PHIC_wea,
        addra     => MPROJ_L1L2G_D3PHIC_writeaddr,
        dina      => MPROJ_L1L2G_D3PHIC_din,
        wea_out       => MPROJ_L1L2G_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D3PHIC_start
      );

    MPROJ_L1L2HI_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D3PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_D3PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_D3PHIC_start,
        nent_o    => MPROJ_L1L2HI_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D3PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D3PHIC_wea,
        addra     => MPROJ_L1L2HI_D3PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_D3PHIC_din,
        wea_out       => MPROJ_L1L2HI_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D3PHIC_start
      );

    MPROJ_L1L2JKL_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D3PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D3PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_D3PHIC_start,
        nent_o    => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D3PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D3PHIC_wea,
        addra     => MPROJ_L1L2JKL_D3PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_D3PHIC_din,
        wea_out       => MPROJ_L1L2JKL_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D3PHIC_start
      );

    MPROJ_L2L3ABCD_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D3PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D3PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D3PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D3PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHIC_wea,
        addra     => MPROJ_L2L3ABCD_D3PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_D3PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_D3PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D3PHIC_start
      );

    MPROJ_D1D2ABCD_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIC_wea_delay,
        addra     => MPROJ_D1D2ABCD_D3PHIC_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D3PHIC_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D3PHIC_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D3PHIC_start,
        nent_o    => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D3PHIC_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHIC_wea,
        addra     => MPROJ_D1D2ABCD_D3PHIC_writeaddr,
        dina      => MPROJ_D1D2ABCD_D3PHIC_din,
        wea_out       => MPROJ_D1D2ABCD_D3PHIC_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D3PHIC_start
      );

    MPROJ_L1D1ABCD_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIC_wea_delay,
        addra     => MPROJ_L1D1ABCD_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D3PHIC_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D3PHIC_start,
        nent_o    => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D3PHIC_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D3PHIC_wea,
        addra     => MPROJ_L1D1ABCD_D3PHIC_writeaddr,
        dina      => MPROJ_L1D1ABCD_D3PHIC_din,
        wea_out       => MPROJ_L1D1ABCD_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D3PHIC_start
      );

    MPROJ_L1D1EFGH_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHIC_wea_delay,
        addra     => MPROJ_L1D1EFGH_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D3PHIC_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D3PHIC_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D3PHIC_start,
        nent_o    => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D3PHIC_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHIC_wea,
        addra     => MPROJ_L1D1EFGH_D3PHIC_writeaddr,
        dina      => MPROJ_L1D1EFGH_D3PHIC_din,
        wea_out       => MPROJ_L1D1EFGH_D3PHIC_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D3PHIC_start
      );

    MPROJ_L2D1ABCD_D3PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIC_wea_delay,
        addra     => MPROJ_L2D1ABCD_D3PHIC_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D3PHIC_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D3PHIC_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D3PHIC_start,
        nent_o    => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D3PHIC_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHIC_wea,
        addra     => MPROJ_L2D1ABCD_D3PHIC_writeaddr,
        dina      => MPROJ_L2D1ABCD_D3PHIC_din,
        wea_out       => MPROJ_L2D1ABCD_D3PHIC_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D3PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D3PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D3PHIC_start
      );

    MPROJ_L1L2G_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D3PHID_wea_delay,
        addra     => MPROJ_L1L2G_D3PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D3PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_D3PHID_V_dout,
        sync_nent => MPROJ_L1L2G_D3PHID_start,
        nent_o    => MPROJ_L1L2G_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D3PHID_AV_dout_mask
      );

    MPROJ_L1L2G_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D3PHID_wea,
        addra     => MPROJ_L1L2G_D3PHID_writeaddr,
        dina      => MPROJ_L1L2G_D3PHID_din,
        wea_out       => MPROJ_L1L2G_D3PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D3PHID_start
      );

    MPROJ_L1L2HI_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D3PHID_wea_delay,
        addra     => MPROJ_L1L2HI_D3PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D3PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_D3PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_D3PHID_start,
        nent_o    => MPROJ_L1L2HI_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D3PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D3PHID_wea,
        addra     => MPROJ_L1L2HI_D3PHID_writeaddr,
        dina      => MPROJ_L1L2HI_D3PHID_din,
        wea_out       => MPROJ_L1L2HI_D3PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D3PHID_start
      );

    MPROJ_L1L2JKL_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D3PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_D3PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D3PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D3PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_D3PHID_start,
        nent_o    => MPROJ_L1L2JKL_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D3PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D3PHID_wea,
        addra     => MPROJ_L1L2JKL_D3PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_D3PHID_din,
        wea_out       => MPROJ_L1L2JKL_D3PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D3PHID_start
      );

    MPROJ_L2L3ABCD_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_D3PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D3PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D3PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D3PHID_start,
        nent_o    => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D3PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D3PHID_wea,
        addra     => MPROJ_L2L3ABCD_D3PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_D3PHID_din,
        wea_out       => MPROJ_L2L3ABCD_D3PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D3PHID_start
      );

    MPROJ_D1D2ABCD_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHID_wea_delay,
        addra     => MPROJ_D1D2ABCD_D3PHID_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D3PHID_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D3PHID_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D3PHID_start,
        nent_o    => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D3PHID_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D3PHID_wea,
        addra     => MPROJ_D1D2ABCD_D3PHID_writeaddr,
        dina      => MPROJ_D1D2ABCD_D3PHID_din,
        wea_out       => MPROJ_D1D2ABCD_D3PHID_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D3PHID_start
      );

    MPROJ_L1D1EFGH_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHID_wea_delay,
        addra     => MPROJ_L1D1EFGH_D3PHID_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D3PHID_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D3PHID_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D3PHID_start,
        nent_o    => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D3PHID_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D3PHID_wea,
        addra     => MPROJ_L1D1EFGH_D3PHID_writeaddr,
        dina      => MPROJ_L1D1EFGH_D3PHID_din,
        wea_out       => MPROJ_L1D1EFGH_D3PHID_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D3PHID_start
      );

    MPROJ_L2D1ABCD_D3PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHID_wea_delay,
        addra     => MPROJ_L2D1ABCD_D3PHID_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D3PHID_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D3PHID_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D3PHID_start,
        nent_o    => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D3PHID_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D3PHID_wea,
        addra     => MPROJ_L2D1ABCD_D3PHID_writeaddr,
        dina      => MPROJ_L2D1ABCD_D3PHID_din,
        wea_out       => MPROJ_L2D1ABCD_D3PHID_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D3PHID_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D3PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D3PHID_start
      );

    MPROJ_L1L2ABC_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D4PHIA_wea_delay,
        addra     => MPROJ_L1L2ABC_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D4PHIA_V_dout,
        sync_nent => MPROJ_L1L2ABC_D4PHIA_start,
        nent_o    => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D4PHIA_AV_dout_mask
      );

    MPROJ_L1L2ABC_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D4PHIA_wea,
        addra     => MPROJ_L1L2ABC_D4PHIA_writeaddr,
        dina      => MPROJ_L1L2ABC_D4PHIA_din,
        wea_out       => MPROJ_L1L2ABC_D4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D4PHIA_start
      );

    MPROJ_L1L2DE_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D4PHIA_wea_delay,
        addra     => MPROJ_L1L2DE_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2DE_D4PHIA_V_dout,
        sync_nent => MPROJ_L1L2DE_D4PHIA_start,
        nent_o    => MPROJ_L1L2DE_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D4PHIA_AV_dout_mask
      );

    MPROJ_L1L2DE_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D4PHIA_wea,
        addra     => MPROJ_L1L2DE_D4PHIA_writeaddr,
        dina      => MPROJ_L1L2DE_D4PHIA_din,
        wea_out       => MPROJ_L1L2DE_D4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2DE_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D4PHIA_start
      );

    MPROJ_L1L2F_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D4PHIA_wea_delay,
        addra     => MPROJ_L1L2F_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L1L2F_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D4PHIA_V_readaddr,
        doutb     => MPROJ_L1L2F_D4PHIA_V_dout,
        sync_nent => MPROJ_L1L2F_D4PHIA_start,
        nent_o    => MPROJ_L1L2F_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D4PHIA_AV_dout_mask
      );

    MPROJ_L1L2F_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D4PHIA_wea,
        addra     => MPROJ_L1L2F_D4PHIA_writeaddr,
        dina      => MPROJ_L1L2F_D4PHIA_din,
        wea_out       => MPROJ_L1L2F_D4PHIA_wea_delay,
        addra_out     => MPROJ_L1L2F_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D4PHIA_start
      );

    MPROJ_L2L3ABCD_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIA_wea_delay,
        addra     => MPROJ_L2L3ABCD_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D4PHIA_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D4PHIA_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D4PHIA_start,
        nent_o    => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D4PHIA_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIA_wea,
        addra     => MPROJ_L2L3ABCD_D4PHIA_writeaddr,
        dina      => MPROJ_L2L3ABCD_D4PHIA_din,
        wea_out       => MPROJ_L2L3ABCD_D4PHIA_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D4PHIA_start
      );

    MPROJ_D1D2ABCD_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIA_wea_delay,
        addra     => MPROJ_D1D2ABCD_D4PHIA_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D4PHIA_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D4PHIA_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D4PHIA_start,
        nent_o    => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D4PHIA_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIA_wea,
        addra     => MPROJ_D1D2ABCD_D4PHIA_writeaddr,
        dina      => MPROJ_D1D2ABCD_D4PHIA_din,
        wea_out       => MPROJ_D1D2ABCD_D4PHIA_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D4PHIA_start
      );

    MPROJ_L1D1ABCD_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIA_wea_delay,
        addra     => MPROJ_L1D1ABCD_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D4PHIA_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D4PHIA_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D4PHIA_start,
        nent_o    => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D4PHIA_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIA_wea,
        addra     => MPROJ_L1D1ABCD_D4PHIA_writeaddr,
        dina      => MPROJ_L1D1ABCD_D4PHIA_din,
        wea_out       => MPROJ_L1D1ABCD_D4PHIA_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D4PHIA_start
      );

    MPROJ_L2D1ABCD_D4PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIA_wea_delay,
        addra     => MPROJ_L2D1ABCD_D4PHIA_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D4PHIA_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D4PHIA_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D4PHIA_start,
        nent_o    => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D4PHIA_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIA_wea,
        addra     => MPROJ_L2D1ABCD_D4PHIA_writeaddr,
        dina      => MPROJ_L2D1ABCD_D4PHIA_din,
        wea_out       => MPROJ_L2D1ABCD_D4PHIA_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D4PHIA_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D4PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D4PHIA_start
      );

    MPROJ_L1L2ABC_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2ABC_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2ABC_D4PHIB_wea_delay,
        addra     => MPROJ_L1L2ABC_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2ABC_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2ABC_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2ABC_D4PHIB_V_dout,
        sync_nent => MPROJ_L1L2ABC_D4PHIB_start,
        nent_o    => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2ABC_D4PHIB_AV_dout_mask
      );

    MPROJ_L1L2ABC_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2ABC_D4PHIB_wea,
        addra     => MPROJ_L1L2ABC_D4PHIB_writeaddr,
        dina      => MPROJ_L1L2ABC_D4PHIB_din,
        wea_out       => MPROJ_L1L2ABC_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2ABC_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2ABC_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2ABC_D4PHIB_start
      );

    MPROJ_L1L2DE_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D4PHIB_wea_delay,
        addra     => MPROJ_L1L2DE_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2DE_D4PHIB_V_dout,
        sync_nent => MPROJ_L1L2DE_D4PHIB_start,
        nent_o    => MPROJ_L1L2DE_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D4PHIB_AV_dout_mask
      );

    MPROJ_L1L2DE_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D4PHIB_wea,
        addra     => MPROJ_L1L2DE_D4PHIB_writeaddr,
        dina      => MPROJ_L1L2DE_D4PHIB_din,
        wea_out       => MPROJ_L1L2DE_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2DE_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D4PHIB_start
      );

    MPROJ_L1L2F_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D4PHIB_wea_delay,
        addra     => MPROJ_L1L2F_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2F_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2F_D4PHIB_V_dout,
        sync_nent => MPROJ_L1L2F_D4PHIB_start,
        nent_o    => MPROJ_L1L2F_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D4PHIB_AV_dout_mask
      );

    MPROJ_L1L2F_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D4PHIB_wea,
        addra     => MPROJ_L1L2F_D4PHIB_writeaddr,
        dina      => MPROJ_L1L2F_D4PHIB_din,
        wea_out       => MPROJ_L1L2F_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2F_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D4PHIB_start
      );

    MPROJ_L1L2G_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D4PHIB_wea_delay,
        addra     => MPROJ_L1L2G_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2G_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2G_D4PHIB_V_dout,
        sync_nent => MPROJ_L1L2G_D4PHIB_start,
        nent_o    => MPROJ_L1L2G_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D4PHIB_AV_dout_mask
      );

    MPROJ_L1L2G_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D4PHIB_wea,
        addra     => MPROJ_L1L2G_D4PHIB_writeaddr,
        dina      => MPROJ_L1L2G_D4PHIB_din,
        wea_out       => MPROJ_L1L2G_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2G_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D4PHIB_start
      );

    MPROJ_L1L2HI_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D4PHIB_wea_delay,
        addra     => MPROJ_L1L2HI_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1L2HI_D4PHIB_V_dout,
        sync_nent => MPROJ_L1L2HI_D4PHIB_start,
        nent_o    => MPROJ_L1L2HI_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D4PHIB_AV_dout_mask
      );

    MPROJ_L1L2HI_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D4PHIB_wea,
        addra     => MPROJ_L1L2HI_D4PHIB_writeaddr,
        dina      => MPROJ_L1L2HI_D4PHIB_din,
        wea_out       => MPROJ_L1L2HI_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1L2HI_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D4PHIB_start
      );

    MPROJ_L2L3ABCD_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIB_wea_delay,
        addra     => MPROJ_L2L3ABCD_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D4PHIB_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D4PHIB_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D4PHIB_start,
        nent_o    => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D4PHIB_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIB_wea,
        addra     => MPROJ_L2L3ABCD_D4PHIB_writeaddr,
        dina      => MPROJ_L2L3ABCD_D4PHIB_din,
        wea_out       => MPROJ_L2L3ABCD_D4PHIB_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D4PHIB_start
      );

    MPROJ_D1D2ABCD_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIB_wea_delay,
        addra     => MPROJ_D1D2ABCD_D4PHIB_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D4PHIB_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D4PHIB_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D4PHIB_start,
        nent_o    => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D4PHIB_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIB_wea,
        addra     => MPROJ_D1D2ABCD_D4PHIB_writeaddr,
        dina      => MPROJ_D1D2ABCD_D4PHIB_din,
        wea_out       => MPROJ_D1D2ABCD_D4PHIB_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D4PHIB_start
      );

    MPROJ_L1D1ABCD_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIB_wea_delay,
        addra     => MPROJ_L1D1ABCD_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D4PHIB_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D4PHIB_start,
        nent_o    => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D4PHIB_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIB_wea,
        addra     => MPROJ_L1D1ABCD_D4PHIB_writeaddr,
        dina      => MPROJ_L1D1ABCD_D4PHIB_din,
        wea_out       => MPROJ_L1D1ABCD_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D4PHIB_start
      );

    MPROJ_L1D1EFGH_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHIB_wea_delay,
        addra     => MPROJ_L1D1EFGH_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D4PHIB_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D4PHIB_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D4PHIB_start,
        nent_o    => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D4PHIB_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHIB_wea,
        addra     => MPROJ_L1D1EFGH_D4PHIB_writeaddr,
        dina      => MPROJ_L1D1EFGH_D4PHIB_din,
        wea_out       => MPROJ_L1D1EFGH_D4PHIB_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D4PHIB_start
      );

    MPROJ_L2D1ABCD_D4PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIB_wea_delay,
        addra     => MPROJ_L2D1ABCD_D4PHIB_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D4PHIB_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D4PHIB_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D4PHIB_start,
        nent_o    => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D4PHIB_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIB_wea,
        addra     => MPROJ_L2D1ABCD_D4PHIB_writeaddr,
        dina      => MPROJ_L2D1ABCD_D4PHIB_din,
        wea_out       => MPROJ_L2D1ABCD_D4PHIB_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D4PHIB_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D4PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D4PHIB_start
      );

    MPROJ_L1L2DE_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2DE_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2DE_D4PHIC_wea_delay,
        addra     => MPROJ_L1L2DE_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2DE_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2DE_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2DE_D4PHIC_V_dout,
        sync_nent => MPROJ_L1L2DE_D4PHIC_start,
        nent_o    => MPROJ_L1L2DE_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2DE_D4PHIC_AV_dout_mask
      );

    MPROJ_L1L2DE_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2DE_D4PHIC_wea,
        addra     => MPROJ_L1L2DE_D4PHIC_writeaddr,
        dina      => MPROJ_L1L2DE_D4PHIC_din,
        wea_out       => MPROJ_L1L2DE_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2DE_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2DE_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2DE_D4PHIC_start
      );

    MPROJ_L1L2F_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2F_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2F_D4PHIC_wea_delay,
        addra     => MPROJ_L1L2F_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2F_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2F_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2F_D4PHIC_V_dout,
        sync_nent => MPROJ_L1L2F_D4PHIC_start,
        nent_o    => MPROJ_L1L2F_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2F_D4PHIC_AV_dout_mask
      );

    MPROJ_L1L2F_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2F_D4PHIC_wea,
        addra     => MPROJ_L1L2F_D4PHIC_writeaddr,
        dina      => MPROJ_L1L2F_D4PHIC_din,
        wea_out       => MPROJ_L1L2F_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2F_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2F_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2F_D4PHIC_start
      );

    MPROJ_L1L2G_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D4PHIC_wea_delay,
        addra     => MPROJ_L1L2G_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2G_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2G_D4PHIC_V_dout,
        sync_nent => MPROJ_L1L2G_D4PHIC_start,
        nent_o    => MPROJ_L1L2G_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D4PHIC_AV_dout_mask
      );

    MPROJ_L1L2G_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D4PHIC_wea,
        addra     => MPROJ_L1L2G_D4PHIC_writeaddr,
        dina      => MPROJ_L1L2G_D4PHIC_din,
        wea_out       => MPROJ_L1L2G_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2G_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D4PHIC_start
      );

    MPROJ_L1L2HI_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D4PHIC_wea_delay,
        addra     => MPROJ_L1L2HI_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2HI_D4PHIC_V_dout,
        sync_nent => MPROJ_L1L2HI_D4PHIC_start,
        nent_o    => MPROJ_L1L2HI_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D4PHIC_AV_dout_mask
      );

    MPROJ_L1L2HI_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D4PHIC_wea,
        addra     => MPROJ_L1L2HI_D4PHIC_writeaddr,
        dina      => MPROJ_L1L2HI_D4PHIC_din,
        wea_out       => MPROJ_L1L2HI_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2HI_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D4PHIC_start
      );

    MPROJ_L1L2JKL_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D4PHIC_wea_delay,
        addra     => MPROJ_L1L2JKL_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D4PHIC_V_dout,
        sync_nent => MPROJ_L1L2JKL_D4PHIC_start,
        nent_o    => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D4PHIC_AV_dout_mask
      );

    MPROJ_L1L2JKL_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D4PHIC_wea,
        addra     => MPROJ_L1L2JKL_D4PHIC_writeaddr,
        dina      => MPROJ_L1L2JKL_D4PHIC_din,
        wea_out       => MPROJ_L1L2JKL_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D4PHIC_start
      );

    MPROJ_L2L3ABCD_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIC_wea_delay,
        addra     => MPROJ_L2L3ABCD_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D4PHIC_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D4PHIC_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D4PHIC_start,
        nent_o    => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D4PHIC_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHIC_wea,
        addra     => MPROJ_L2L3ABCD_D4PHIC_writeaddr,
        dina      => MPROJ_L2L3ABCD_D4PHIC_din,
        wea_out       => MPROJ_L2L3ABCD_D4PHIC_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D4PHIC_start
      );

    MPROJ_D1D2ABCD_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIC_wea_delay,
        addra     => MPROJ_D1D2ABCD_D4PHIC_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D4PHIC_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D4PHIC_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D4PHIC_start,
        nent_o    => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D4PHIC_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHIC_wea,
        addra     => MPROJ_D1D2ABCD_D4PHIC_writeaddr,
        dina      => MPROJ_D1D2ABCD_D4PHIC_din,
        wea_out       => MPROJ_D1D2ABCD_D4PHIC_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D4PHIC_start
      );

    MPROJ_L1D1ABCD_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIC_wea_delay,
        addra     => MPROJ_L1D1ABCD_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D4PHIC_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D4PHIC_start,
        nent_o    => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D4PHIC_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D4PHIC_wea,
        addra     => MPROJ_L1D1ABCD_D4PHIC_writeaddr,
        dina      => MPROJ_L1D1ABCD_D4PHIC_din,
        wea_out       => MPROJ_L1D1ABCD_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D4PHIC_start
      );

    MPROJ_L1D1EFGH_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHIC_wea_delay,
        addra     => MPROJ_L1D1EFGH_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D4PHIC_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D4PHIC_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D4PHIC_start,
        nent_o    => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D4PHIC_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHIC_wea,
        addra     => MPROJ_L1D1EFGH_D4PHIC_writeaddr,
        dina      => MPROJ_L1D1EFGH_D4PHIC_din,
        wea_out       => MPROJ_L1D1EFGH_D4PHIC_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D4PHIC_start
      );

    MPROJ_L2D1ABCD_D4PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIC_wea_delay,
        addra     => MPROJ_L2D1ABCD_D4PHIC_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D4PHIC_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D4PHIC_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D4PHIC_start,
        nent_o    => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D4PHIC_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHIC_wea,
        addra     => MPROJ_L2D1ABCD_D4PHIC_writeaddr,
        dina      => MPROJ_L2D1ABCD_D4PHIC_din,
        wea_out       => MPROJ_L2D1ABCD_D4PHIC_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D4PHIC_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D4PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D4PHIC_start
      );

    MPROJ_L1L2G_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2G_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2G_D4PHID_wea_delay,
        addra     => MPROJ_L1L2G_D4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2G_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2G_D4PHID_V_readaddr,
        doutb     => MPROJ_L1L2G_D4PHID_V_dout,
        sync_nent => MPROJ_L1L2G_D4PHID_start,
        nent_o    => MPROJ_L1L2G_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2G_D4PHID_AV_dout_mask
      );

    MPROJ_L1L2G_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2G_D4PHID_wea,
        addra     => MPROJ_L1L2G_D4PHID_writeaddr,
        dina      => MPROJ_L1L2G_D4PHID_din,
        wea_out       => MPROJ_L1L2G_D4PHID_wea_delay,
        addra_out     => MPROJ_L1L2G_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2G_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2G_D4PHID_start
      );

    MPROJ_L1L2HI_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2HI_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2HI_D4PHID_wea_delay,
        addra     => MPROJ_L1L2HI_D4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2HI_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2HI_D4PHID_V_readaddr,
        doutb     => MPROJ_L1L2HI_D4PHID_V_dout,
        sync_nent => MPROJ_L1L2HI_D4PHID_start,
        nent_o    => MPROJ_L1L2HI_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2HI_D4PHID_AV_dout_mask
      );

    MPROJ_L1L2HI_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2HI_D4PHID_wea,
        addra     => MPROJ_L1L2HI_D4PHID_writeaddr,
        dina      => MPROJ_L1L2HI_D4PHID_din,
        wea_out       => MPROJ_L1L2HI_D4PHID_wea_delay,
        addra_out     => MPROJ_L1L2HI_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2HI_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2HI_D4PHID_start
      );

    MPROJ_L1L2JKL_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1L2JKL_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1L2JKL_D4PHID_wea_delay,
        addra     => MPROJ_L1L2JKL_D4PHID_writeaddr_delay,
        dina      => MPROJ_L1L2JKL_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1L2JKL_D4PHID_V_readaddr,
        doutb     => MPROJ_L1L2JKL_D4PHID_V_dout,
        sync_nent => MPROJ_L1L2JKL_D4PHID_start,
        nent_o    => MPROJ_L1L2JKL_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1L2JKL_D4PHID_AV_dout_mask
      );

    MPROJ_L1L2JKL_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1L2JKL_D4PHID_wea,
        addra     => MPROJ_L1L2JKL_D4PHID_writeaddr,
        dina      => MPROJ_L1L2JKL_D4PHID_din,
        wea_out       => MPROJ_L1L2JKL_D4PHID_wea_delay,
        addra_out     => MPROJ_L1L2JKL_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1L2JKL_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1L2JKL_D4PHID_start
      );

    MPROJ_L2L3ABCD_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2L3ABCD_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHID_wea_delay,
        addra     => MPROJ_L2L3ABCD_D4PHID_writeaddr_delay,
        dina      => MPROJ_L2L3ABCD_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2L3ABCD_D4PHID_V_readaddr,
        doutb     => MPROJ_L2L3ABCD_D4PHID_V_dout,
        sync_nent => MPROJ_L2L3ABCD_D4PHID_start,
        nent_o    => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L2L3ABCD_D4PHID_AV_dout_mask
      );

    MPROJ_L2L3ABCD_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2L3ABCD_D4PHID_wea,
        addra     => MPROJ_L2L3ABCD_D4PHID_writeaddr,
        dina      => MPROJ_L2L3ABCD_D4PHID_din,
        wea_out       => MPROJ_L2L3ABCD_D4PHID_wea_delay,
        addra_out     => MPROJ_L2L3ABCD_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L2L3ABCD_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2L3ABCD_D4PHID_start
      );

    MPROJ_D1D2ABCD_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHID_wea_delay,
        addra     => MPROJ_D1D2ABCD_D4PHID_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D4PHID_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D4PHID_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D4PHID_start,
        nent_o    => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D4PHID_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D4PHID_wea,
        addra     => MPROJ_D1D2ABCD_D4PHID_writeaddr,
        dina      => MPROJ_D1D2ABCD_D4PHID_din,
        wea_out       => MPROJ_D1D2ABCD_D4PHID_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D4PHID_start
      );

    MPROJ_L1D1EFGH_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHID_wea_delay,
        addra     => MPROJ_L1D1EFGH_D4PHID_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D4PHID_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D4PHID_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D4PHID_start,
        nent_o    => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D4PHID_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D4PHID_wea,
        addra     => MPROJ_L1D1EFGH_D4PHID_writeaddr,
        dina      => MPROJ_L1D1EFGH_D4PHID_din,
        wea_out       => MPROJ_L1D1EFGH_D4PHID_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D4PHID_start
      );

    MPROJ_L2D1ABCD_D4PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L2D1ABCD_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHID_wea_delay,
        addra     => MPROJ_L2D1ABCD_D4PHID_writeaddr_delay,
        dina      => MPROJ_L2D1ABCD_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L2D1ABCD_D4PHID_V_readaddr,
        doutb     => MPROJ_L2D1ABCD_D4PHID_V_dout,
        sync_nent => MPROJ_L2D1ABCD_D4PHID_start,
        nent_o    => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent,
        mask_o    => MPROJ_L2D1ABCD_D4PHID_AV_dout_mask
      );

    MPROJ_L2D1ABCD_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L2D1ABCD_D4PHID_wea,
        addra     => MPROJ_L2D1ABCD_D4PHID_writeaddr,
        dina      => MPROJ_L2D1ABCD_D4PHID_din,
        wea_out       => MPROJ_L2D1ABCD_D4PHID_wea_delay,
        addra_out     => MPROJ_L2D1ABCD_D4PHID_writeaddr_delay,
        dina_out      => MPROJ_L2D1ABCD_D4PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L2D1ABCD_D4PHID_start
      );

    MPROJ_D1D2ABCD_D5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIA_wea_delay,
        addra     => MPROJ_D1D2ABCD_D5PHIA_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D5PHIA_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D5PHIA_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D5PHIA_start,
        nent_o    => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D5PHIA_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIA_wea,
        addra     => MPROJ_D1D2ABCD_D5PHIA_writeaddr,
        dina      => MPROJ_D1D2ABCD_D5PHIA_din,
        wea_out       => MPROJ_D1D2ABCD_D5PHIA_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D5PHIA_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D5PHIA_start
      );

    MPROJ_D3D4ABCD_D5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIA_wea_delay,
        addra     => MPROJ_D3D4ABCD_D5PHIA_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D5PHIA_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D5PHIA_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D5PHIA_start,
        nent_o    => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D5PHIA_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIA_wea,
        addra     => MPROJ_D3D4ABCD_D5PHIA_writeaddr,
        dina      => MPROJ_D3D4ABCD_D5PHIA_din,
        wea_out       => MPROJ_D3D4ABCD_D5PHIA_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D5PHIA_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D5PHIA_start
      );

    MPROJ_L1D1ABCD_D5PHIA : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D5PHIA"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIA_wea_delay,
        addra     => MPROJ_L1D1ABCD_D5PHIA_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D5PHIA_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D5PHIA_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D5PHIA_start,
        nent_o    => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D5PHIA_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIA_wea,
        addra     => MPROJ_L1D1ABCD_D5PHIA_writeaddr,
        dina      => MPROJ_L1D1ABCD_D5PHIA_din,
        wea_out       => MPROJ_L1D1ABCD_D5PHIA_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D5PHIA_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D5PHIA_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D5PHIA_start
      );

    MPROJ_D1D2ABCD_D5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIB_wea_delay,
        addra     => MPROJ_D1D2ABCD_D5PHIB_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D5PHIB_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D5PHIB_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D5PHIB_start,
        nent_o    => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D5PHIB_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIB_wea,
        addra     => MPROJ_D1D2ABCD_D5PHIB_writeaddr,
        dina      => MPROJ_D1D2ABCD_D5PHIB_din,
        wea_out       => MPROJ_D1D2ABCD_D5PHIB_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D5PHIB_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D5PHIB_start
      );

    MPROJ_D3D4ABCD_D5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIB_wea_delay,
        addra     => MPROJ_D3D4ABCD_D5PHIB_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D5PHIB_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D5PHIB_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D5PHIB_start,
        nent_o    => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D5PHIB_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIB_wea,
        addra     => MPROJ_D3D4ABCD_D5PHIB_writeaddr,
        dina      => MPROJ_D3D4ABCD_D5PHIB_din,
        wea_out       => MPROJ_D3D4ABCD_D5PHIB_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D5PHIB_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D5PHIB_start
      );

    MPROJ_L1D1ABCD_D5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIB_wea_delay,
        addra     => MPROJ_L1D1ABCD_D5PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D5PHIB_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D5PHIB_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D5PHIB_start,
        nent_o    => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D5PHIB_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIB_wea,
        addra     => MPROJ_L1D1ABCD_D5PHIB_writeaddr,
        dina      => MPROJ_L1D1ABCD_D5PHIB_din,
        wea_out       => MPROJ_L1D1ABCD_D5PHIB_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D5PHIB_start
      );

    MPROJ_L1D1EFGH_D5PHIB : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHIB_wea_delay,
        addra     => MPROJ_L1D1EFGH_D5PHIB_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D5PHIB_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D5PHIB_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D5PHIB_start,
        nent_o    => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D5PHIB_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHIB_wea,
        addra     => MPROJ_L1D1EFGH_D5PHIB_writeaddr,
        dina      => MPROJ_L1D1EFGH_D5PHIB_din,
        wea_out       => MPROJ_L1D1EFGH_D5PHIB_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D5PHIB_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D5PHIB_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D5PHIB_start
      );

    MPROJ_D1D2ABCD_D5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIC_wea_delay,
        addra     => MPROJ_D1D2ABCD_D5PHIC_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D5PHIC_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D5PHIC_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D5PHIC_start,
        nent_o    => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D5PHIC_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHIC_wea,
        addra     => MPROJ_D1D2ABCD_D5PHIC_writeaddr,
        dina      => MPROJ_D1D2ABCD_D5PHIC_din,
        wea_out       => MPROJ_D1D2ABCD_D5PHIC_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D5PHIC_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D5PHIC_start
      );

    MPROJ_D3D4ABCD_D5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIC_wea_delay,
        addra     => MPROJ_D3D4ABCD_D5PHIC_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D5PHIC_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D5PHIC_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D5PHIC_start,
        nent_o    => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D5PHIC_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHIC_wea,
        addra     => MPROJ_D3D4ABCD_D5PHIC_writeaddr,
        dina      => MPROJ_D3D4ABCD_D5PHIC_din,
        wea_out       => MPROJ_D3D4ABCD_D5PHIC_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D5PHIC_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D5PHIC_start
      );

    MPROJ_L1D1ABCD_D5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1ABCD_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIC_wea_delay,
        addra     => MPROJ_L1D1ABCD_D5PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1ABCD_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1ABCD_D5PHIC_V_readaddr,
        doutb     => MPROJ_L1D1ABCD_D5PHIC_V_dout,
        sync_nent => MPROJ_L1D1ABCD_D5PHIC_start,
        nent_o    => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1ABCD_D5PHIC_AV_dout_mask
      );

    MPROJ_L1D1ABCD_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1ABCD_D5PHIC_wea,
        addra     => MPROJ_L1D1ABCD_D5PHIC_writeaddr,
        dina      => MPROJ_L1D1ABCD_D5PHIC_din,
        wea_out       => MPROJ_L1D1ABCD_D5PHIC_wea_delay,
        addra_out     => MPROJ_L1D1ABCD_D5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1ABCD_D5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1ABCD_D5PHIC_start
      );

    MPROJ_L1D1EFGH_D5PHIC : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHIC_wea_delay,
        addra     => MPROJ_L1D1EFGH_D5PHIC_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D5PHIC_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D5PHIC_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D5PHIC_start,
        nent_o    => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D5PHIC_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHIC_wea,
        addra     => MPROJ_L1D1EFGH_D5PHIC_writeaddr,
        dina      => MPROJ_L1D1EFGH_D5PHIC_din,
        wea_out       => MPROJ_L1D1EFGH_D5PHIC_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D5PHIC_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D5PHIC_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D5PHIC_start
      );

    MPROJ_D1D2ABCD_D5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D1D2ABCD_D5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHID_wea_delay,
        addra     => MPROJ_D1D2ABCD_D5PHID_writeaddr_delay,
        dina      => MPROJ_D1D2ABCD_D5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D1D2ABCD_D5PHID_V_readaddr,
        doutb     => MPROJ_D1D2ABCD_D5PHID_V_dout,
        sync_nent => MPROJ_D1D2ABCD_D5PHID_start,
        nent_o    => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent,
        mask_o    => MPROJ_D1D2ABCD_D5PHID_AV_dout_mask
      );

    MPROJ_D1D2ABCD_D5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D1D2ABCD_D5PHID_wea,
        addra     => MPROJ_D1D2ABCD_D5PHID_writeaddr,
        dina      => MPROJ_D1D2ABCD_D5PHID_din,
        wea_out       => MPROJ_D1D2ABCD_D5PHID_wea_delay,
        addra_out     => MPROJ_D1D2ABCD_D5PHID_writeaddr_delay,
        dina_out      => MPROJ_D1D2ABCD_D5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D1D2ABCD_D5PHID_start
      );

    MPROJ_D3D4ABCD_D5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_D3D4ABCD_D5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHID_wea_delay,
        addra     => MPROJ_D3D4ABCD_D5PHID_writeaddr_delay,
        dina      => MPROJ_D3D4ABCD_D5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_D3D4ABCD_D5PHID_V_readaddr,
        doutb     => MPROJ_D3D4ABCD_D5PHID_V_dout,
        sync_nent => MPROJ_D3D4ABCD_D5PHID_start,
        nent_o    => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent,
        mask_o    => MPROJ_D3D4ABCD_D5PHID_AV_dout_mask
      );

    MPROJ_D3D4ABCD_D5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_D3D4ABCD_D5PHID_wea,
        addra     => MPROJ_D3D4ABCD_D5PHID_writeaddr,
        dina      => MPROJ_D3D4ABCD_D5PHID_din,
        wea_out       => MPROJ_D3D4ABCD_D5PHID_wea_delay,
        addra_out     => MPROJ_D3D4ABCD_D5PHID_writeaddr_delay,
        dina_out      => MPROJ_D3D4ABCD_D5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_D3D4ABCD_D5PHID_start
      );

    MPROJ_L1D1EFGH_D5PHID : entity work.tf_mem_tproj
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        PAGE_LENGTH       => 64,
        NUM_TPAGES       => 4,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "MPROJ_L1D1EFGH_D5PHID"
      )
      port map (
        clka      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHID_wea_delay,
        addra     => MPROJ_L1D1EFGH_D5PHID_writeaddr_delay,
        dina      => MPROJ_L1D1EFGH_D5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => MPROJ_L1D1EFGH_D5PHID_V_readaddr,
        doutb     => MPROJ_L1D1EFGH_D5PHID_V_dout,
        sync_nent => MPROJ_L1D1EFGH_D5PHID_start,
        nent_o    => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent,
        mask_o    => MPROJ_L1D1EFGH_D5PHID_AV_dout_mask
      );

    MPROJ_L1D1EFGH_D5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        PAGE_LENGTH       => 64,
        NUM_PAGES       => 8,
        RAM_WIDTH       => 59
      )
      port map (
        clk      => clk,
        wea       => MPROJ_L1D1EFGH_D5PHID_wea,
        addra     => MPROJ_L1D1EFGH_D5PHID_writeaddr,
        dina      => MPROJ_L1D1EFGH_D5PHID_din,
        wea_out       => MPROJ_L1D1EFGH_D5PHID_wea_delay,
        addra_out     => MPROJ_L1D1EFGH_D5PHID_writeaddr_delay,
        dina_out      => MPROJ_L1D1EFGH_D5PHID_din_delay,
        done       => PC_done,
        start      => MPROJ_L1D1EFGH_D5PHID_start
      );

    FM_AAAA_L1PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIA_wea_delay,
        addra     => FM_AAAA_L1PHIA_writeaddr_delay,
        dina      => FM_AAAA_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIA_V_readaddr,
        doutb     => FM_AAAA_L1PHIA_V_dout,
        sync_nent => FM_AAAA_L1PHIA_start,
        nent_o    => FM_AAAA_L1PHIA_AV_dout_nent
      );

    FM_AAAA_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIA_wea,
        addra     => FM_AAAA_L1PHIA_writeaddr,
        dina      => FM_AAAA_L1PHIA_din,
        wea_out       => FM_AAAA_L1PHIA_wea_delay,
        addra_out     => FM_AAAA_L1PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIA_start
      );

    FM_BBBB_L1PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIA_wea_delay,
        addra     => FM_BBBB_L1PHIA_writeaddr_delay,
        dina      => FM_BBBB_L1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIA_V_readaddr,
        doutb     => FM_BBBB_L1PHIA_V_dout,
        sync_nent => FM_BBBB_L1PHIA_start,
        nent_o    => FM_BBBB_L1PHIA_AV_dout_nent
      );

    FM_BBBB_L1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIA_wea,
        addra     => FM_BBBB_L1PHIA_writeaddr,
        dina      => FM_BBBB_L1PHIA_din,
        wea_out       => FM_BBBB_L1PHIA_wea_delay,
        addra_out     => FM_BBBB_L1PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIA_start
      );

    FM_AAAA_L1PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIB_wea_delay,
        addra     => FM_AAAA_L1PHIB_writeaddr_delay,
        dina      => FM_AAAA_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIB_V_readaddr,
        doutb     => FM_AAAA_L1PHIB_V_dout,
        sync_nent => FM_AAAA_L1PHIB_start,
        nent_o    => FM_AAAA_L1PHIB_AV_dout_nent
      );

    FM_AAAA_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIB_wea,
        addra     => FM_AAAA_L1PHIB_writeaddr,
        dina      => FM_AAAA_L1PHIB_din,
        wea_out       => FM_AAAA_L1PHIB_wea_delay,
        addra_out     => FM_AAAA_L1PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIB_start
      );

    FM_BBBB_L1PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIB_wea_delay,
        addra     => FM_BBBB_L1PHIB_writeaddr_delay,
        dina      => FM_BBBB_L1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIB_V_readaddr,
        doutb     => FM_BBBB_L1PHIB_V_dout,
        sync_nent => FM_BBBB_L1PHIB_start,
        nent_o    => FM_BBBB_L1PHIB_AV_dout_nent
      );

    FM_BBBB_L1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIB_wea,
        addra     => FM_BBBB_L1PHIB_writeaddr,
        dina      => FM_BBBB_L1PHIB_din,
        wea_out       => FM_BBBB_L1PHIB_wea_delay,
        addra_out     => FM_BBBB_L1PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIB_start
      );

    FM_AAAA_L1PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIC_wea_delay,
        addra     => FM_AAAA_L1PHIC_writeaddr_delay,
        dina      => FM_AAAA_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIC_V_readaddr,
        doutb     => FM_AAAA_L1PHIC_V_dout,
        sync_nent => FM_AAAA_L1PHIC_start,
        nent_o    => FM_AAAA_L1PHIC_AV_dout_nent
      );

    FM_AAAA_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIC_wea,
        addra     => FM_AAAA_L1PHIC_writeaddr,
        dina      => FM_AAAA_L1PHIC_din,
        wea_out       => FM_AAAA_L1PHIC_wea_delay,
        addra_out     => FM_AAAA_L1PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIC_start
      );

    FM_BBBB_L1PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIC_wea_delay,
        addra     => FM_BBBB_L1PHIC_writeaddr_delay,
        dina      => FM_BBBB_L1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIC_V_readaddr,
        doutb     => FM_BBBB_L1PHIC_V_dout,
        sync_nent => FM_BBBB_L1PHIC_start,
        nent_o    => FM_BBBB_L1PHIC_AV_dout_nent
      );

    FM_BBBB_L1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIC_wea,
        addra     => FM_BBBB_L1PHIC_writeaddr,
        dina      => FM_BBBB_L1PHIC_din,
        wea_out       => FM_BBBB_L1PHIC_wea_delay,
        addra_out     => FM_BBBB_L1PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIC_start
      );

    FM_AAAA_L1PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHID_wea_delay,
        addra     => FM_AAAA_L1PHID_writeaddr_delay,
        dina      => FM_AAAA_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHID_V_readaddr,
        doutb     => FM_AAAA_L1PHID_V_dout,
        sync_nent => FM_AAAA_L1PHID_start,
        nent_o    => FM_AAAA_L1PHID_AV_dout_nent
      );

    FM_AAAA_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHID_wea,
        addra     => FM_AAAA_L1PHID_writeaddr,
        dina      => FM_AAAA_L1PHID_din,
        wea_out       => FM_AAAA_L1PHID_wea_delay,
        addra_out     => FM_AAAA_L1PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHID_start
      );

    FM_BBBB_L1PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHID_wea_delay,
        addra     => FM_BBBB_L1PHID_writeaddr_delay,
        dina      => FM_BBBB_L1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHID_V_readaddr,
        doutb     => FM_BBBB_L1PHID_V_dout,
        sync_nent => FM_BBBB_L1PHID_start,
        nent_o    => FM_BBBB_L1PHID_AV_dout_nent
      );

    FM_BBBB_L1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHID_wea,
        addra     => FM_BBBB_L1PHID_writeaddr,
        dina      => FM_BBBB_L1PHID_din,
        wea_out       => FM_BBBB_L1PHID_wea_delay,
        addra_out     => FM_BBBB_L1PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHID_start
      );

    FM_AAAA_L1PHIE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIE_wea_delay,
        addra     => FM_AAAA_L1PHIE_writeaddr_delay,
        dina      => FM_AAAA_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIE_V_readaddr,
        doutb     => FM_AAAA_L1PHIE_V_dout,
        sync_nent => FM_AAAA_L1PHIE_start,
        nent_o    => FM_AAAA_L1PHIE_AV_dout_nent
      );

    FM_AAAA_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIE_wea,
        addra     => FM_AAAA_L1PHIE_writeaddr,
        dina      => FM_AAAA_L1PHIE_din,
        wea_out       => FM_AAAA_L1PHIE_wea_delay,
        addra_out     => FM_AAAA_L1PHIE_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIE_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIE_start
      );

    FM_BBBB_L1PHIE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIE"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIE_wea_delay,
        addra     => FM_BBBB_L1PHIE_writeaddr_delay,
        dina      => FM_BBBB_L1PHIE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIE_V_readaddr,
        doutb     => FM_BBBB_L1PHIE_V_dout,
        sync_nent => FM_BBBB_L1PHIE_start,
        nent_o    => FM_BBBB_L1PHIE_AV_dout_nent
      );

    FM_BBBB_L1PHIE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIE_wea,
        addra     => FM_BBBB_L1PHIE_writeaddr,
        dina      => FM_BBBB_L1PHIE_din,
        wea_out       => FM_BBBB_L1PHIE_wea_delay,
        addra_out     => FM_BBBB_L1PHIE_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIE_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIE_start
      );

    FM_AAAA_L1PHIF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIF_wea_delay,
        addra     => FM_AAAA_L1PHIF_writeaddr_delay,
        dina      => FM_AAAA_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIF_V_readaddr,
        doutb     => FM_AAAA_L1PHIF_V_dout,
        sync_nent => FM_AAAA_L1PHIF_start,
        nent_o    => FM_AAAA_L1PHIF_AV_dout_nent
      );

    FM_AAAA_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIF_wea,
        addra     => FM_AAAA_L1PHIF_writeaddr,
        dina      => FM_AAAA_L1PHIF_din,
        wea_out       => FM_AAAA_L1PHIF_wea_delay,
        addra_out     => FM_AAAA_L1PHIF_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIF_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIF_start
      );

    FM_BBBB_L1PHIF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIF"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIF_wea_delay,
        addra     => FM_BBBB_L1PHIF_writeaddr_delay,
        dina      => FM_BBBB_L1PHIF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIF_V_readaddr,
        doutb     => FM_BBBB_L1PHIF_V_dout,
        sync_nent => FM_BBBB_L1PHIF_start,
        nent_o    => FM_BBBB_L1PHIF_AV_dout_nent
      );

    FM_BBBB_L1PHIF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIF_wea,
        addra     => FM_BBBB_L1PHIF_writeaddr,
        dina      => FM_BBBB_L1PHIF_din,
        wea_out       => FM_BBBB_L1PHIF_wea_delay,
        addra_out     => FM_BBBB_L1PHIF_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIF_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIF_start
      );

    FM_AAAA_L1PHIG : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIG_wea_delay,
        addra     => FM_AAAA_L1PHIG_writeaddr_delay,
        dina      => FM_AAAA_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIG_V_readaddr,
        doutb     => FM_AAAA_L1PHIG_V_dout,
        sync_nent => FM_AAAA_L1PHIG_start,
        nent_o    => FM_AAAA_L1PHIG_AV_dout_nent
      );

    FM_AAAA_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIG_wea,
        addra     => FM_AAAA_L1PHIG_writeaddr,
        dina      => FM_AAAA_L1PHIG_din,
        wea_out       => FM_AAAA_L1PHIG_wea_delay,
        addra_out     => FM_AAAA_L1PHIG_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIG_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIG_start
      );

    FM_BBBB_L1PHIG : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIG"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIG_wea_delay,
        addra     => FM_BBBB_L1PHIG_writeaddr_delay,
        dina      => FM_BBBB_L1PHIG_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIG_V_readaddr,
        doutb     => FM_BBBB_L1PHIG_V_dout,
        sync_nent => FM_BBBB_L1PHIG_start,
        nent_o    => FM_BBBB_L1PHIG_AV_dout_nent
      );

    FM_BBBB_L1PHIG_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIG_wea,
        addra     => FM_BBBB_L1PHIG_writeaddr,
        dina      => FM_BBBB_L1PHIG_din,
        wea_out       => FM_BBBB_L1PHIG_wea_delay,
        addra_out     => FM_BBBB_L1PHIG_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIG_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIG_start
      );

    FM_AAAA_L1PHIH : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L1PHIH_wea_delay,
        addra     => FM_AAAA_L1PHIH_writeaddr_delay,
        dina      => FM_AAAA_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L1PHIH_V_readaddr,
        doutb     => FM_AAAA_L1PHIH_V_dout,
        sync_nent => FM_AAAA_L1PHIH_start,
        nent_o    => FM_AAAA_L1PHIH_AV_dout_nent
      );

    FM_AAAA_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L1PHIH_wea,
        addra     => FM_AAAA_L1PHIH_writeaddr,
        dina      => FM_AAAA_L1PHIH_din,
        wea_out       => FM_AAAA_L1PHIH_wea_delay,
        addra_out     => FM_AAAA_L1PHIH_writeaddr_delay,
        dina_out      => FM_AAAA_L1PHIH_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L1PHIH_start
      );

    FM_BBBB_L1PHIH : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L1PHIH"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L1PHIH_wea_delay,
        addra     => FM_BBBB_L1PHIH_writeaddr_delay,
        dina      => FM_BBBB_L1PHIH_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L1PHIH_V_readaddr,
        doutb     => FM_BBBB_L1PHIH_V_dout,
        sync_nent => FM_BBBB_L1PHIH_start,
        nent_o    => FM_BBBB_L1PHIH_AV_dout_nent
      );

    FM_BBBB_L1PHIH_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L1PHIH_wea,
        addra     => FM_BBBB_L1PHIH_writeaddr,
        dina      => FM_BBBB_L1PHIH_din,
        wea_out       => FM_BBBB_L1PHIH_wea_delay,
        addra_out     => FM_BBBB_L1PHIH_writeaddr_delay,
        dina_out      => FM_BBBB_L1PHIH_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L1PHIH_start
      );

    FM_AAAA_L2PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L2PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L2PHIA_wea_delay,
        addra     => FM_AAAA_L2PHIA_writeaddr_delay,
        dina      => FM_AAAA_L2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L2PHIA_V_readaddr,
        doutb     => FM_AAAA_L2PHIA_V_dout,
        sync_nent => FM_AAAA_L2PHIA_start,
        nent_o    => FM_AAAA_L2PHIA_AV_dout_nent
      );

    FM_AAAA_L2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L2PHIA_wea,
        addra     => FM_AAAA_L2PHIA_writeaddr,
        dina      => FM_AAAA_L2PHIA_din,
        wea_out       => FM_AAAA_L2PHIA_wea_delay,
        addra_out     => FM_AAAA_L2PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L2PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L2PHIA_start
      );

    FM_BBBB_L2PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L2PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L2PHIA_wea_delay,
        addra     => FM_BBBB_L2PHIA_writeaddr_delay,
        dina      => FM_BBBB_L2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L2PHIA_V_readaddr,
        doutb     => FM_BBBB_L2PHIA_V_dout,
        sync_nent => FM_BBBB_L2PHIA_start,
        nent_o    => FM_BBBB_L2PHIA_AV_dout_nent
      );

    FM_BBBB_L2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L2PHIA_wea,
        addra     => FM_BBBB_L2PHIA_writeaddr,
        dina      => FM_BBBB_L2PHIA_din,
        wea_out       => FM_BBBB_L2PHIA_wea_delay,
        addra_out     => FM_BBBB_L2PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L2PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L2PHIA_start
      );

    FM_AAAA_L2PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L2PHIB_wea_delay,
        addra     => FM_AAAA_L2PHIB_writeaddr_delay,
        dina      => FM_AAAA_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L2PHIB_V_readaddr,
        doutb     => FM_AAAA_L2PHIB_V_dout,
        sync_nent => FM_AAAA_L2PHIB_start,
        nent_o    => FM_AAAA_L2PHIB_AV_dout_nent
      );

    FM_AAAA_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L2PHIB_wea,
        addra     => FM_AAAA_L2PHIB_writeaddr,
        dina      => FM_AAAA_L2PHIB_din,
        wea_out       => FM_AAAA_L2PHIB_wea_delay,
        addra_out     => FM_AAAA_L2PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L2PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L2PHIB_start
      );

    FM_BBBB_L2PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L2PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L2PHIB_wea_delay,
        addra     => FM_BBBB_L2PHIB_writeaddr_delay,
        dina      => FM_BBBB_L2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L2PHIB_V_readaddr,
        doutb     => FM_BBBB_L2PHIB_V_dout,
        sync_nent => FM_BBBB_L2PHIB_start,
        nent_o    => FM_BBBB_L2PHIB_AV_dout_nent
      );

    FM_BBBB_L2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L2PHIB_wea,
        addra     => FM_BBBB_L2PHIB_writeaddr,
        dina      => FM_BBBB_L2PHIB_din,
        wea_out       => FM_BBBB_L2PHIB_wea_delay,
        addra_out     => FM_BBBB_L2PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L2PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L2PHIB_start
      );

    FM_AAAA_L2PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L2PHIC_wea_delay,
        addra     => FM_AAAA_L2PHIC_writeaddr_delay,
        dina      => FM_AAAA_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L2PHIC_V_readaddr,
        doutb     => FM_AAAA_L2PHIC_V_dout,
        sync_nent => FM_AAAA_L2PHIC_start,
        nent_o    => FM_AAAA_L2PHIC_AV_dout_nent
      );

    FM_AAAA_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L2PHIC_wea,
        addra     => FM_AAAA_L2PHIC_writeaddr,
        dina      => FM_AAAA_L2PHIC_din,
        wea_out       => FM_AAAA_L2PHIC_wea_delay,
        addra_out     => FM_AAAA_L2PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L2PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L2PHIC_start
      );

    FM_BBBB_L2PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L2PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L2PHIC_wea_delay,
        addra     => FM_BBBB_L2PHIC_writeaddr_delay,
        dina      => FM_BBBB_L2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L2PHIC_V_readaddr,
        doutb     => FM_BBBB_L2PHIC_V_dout,
        sync_nent => FM_BBBB_L2PHIC_start,
        nent_o    => FM_BBBB_L2PHIC_AV_dout_nent
      );

    FM_BBBB_L2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L2PHIC_wea,
        addra     => FM_BBBB_L2PHIC_writeaddr,
        dina      => FM_BBBB_L2PHIC_din,
        wea_out       => FM_BBBB_L2PHIC_wea_delay,
        addra_out     => FM_BBBB_L2PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L2PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L2PHIC_start
      );

    FM_AAAA_L2PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L2PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L2PHID_wea_delay,
        addra     => FM_AAAA_L2PHID_writeaddr_delay,
        dina      => FM_AAAA_L2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L2PHID_V_readaddr,
        doutb     => FM_AAAA_L2PHID_V_dout,
        sync_nent => FM_AAAA_L2PHID_start,
        nent_o    => FM_AAAA_L2PHID_AV_dout_nent
      );

    FM_AAAA_L2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L2PHID_wea,
        addra     => FM_AAAA_L2PHID_writeaddr,
        dina      => FM_AAAA_L2PHID_din,
        wea_out       => FM_AAAA_L2PHID_wea_delay,
        addra_out     => FM_AAAA_L2PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L2PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L2PHID_start
      );

    FM_BBBB_L2PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L2PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L2PHID_wea_delay,
        addra     => FM_BBBB_L2PHID_writeaddr_delay,
        dina      => FM_BBBB_L2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L2PHID_V_readaddr,
        doutb     => FM_BBBB_L2PHID_V_dout,
        sync_nent => FM_BBBB_L2PHID_start,
        nent_o    => FM_BBBB_L2PHID_AV_dout_nent
      );

    FM_BBBB_L2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L2PHID_wea,
        addra     => FM_BBBB_L2PHID_writeaddr,
        dina      => FM_BBBB_L2PHID_din,
        wea_out       => FM_BBBB_L2PHID_wea_delay,
        addra_out     => FM_BBBB_L2PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L2PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L2PHID_start
      );

    FM_AAAA_L3PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L3PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L3PHIA_wea_delay,
        addra     => FM_AAAA_L3PHIA_writeaddr_delay,
        dina      => FM_AAAA_L3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L3PHIA_V_readaddr,
        doutb     => FM_AAAA_L3PHIA_V_dout,
        sync_nent => FM_AAAA_L3PHIA_start,
        nent_o    => FM_AAAA_L3PHIA_AV_dout_nent
      );

    FM_AAAA_L3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L3PHIA_wea,
        addra     => FM_AAAA_L3PHIA_writeaddr,
        dina      => FM_AAAA_L3PHIA_din,
        wea_out       => FM_AAAA_L3PHIA_wea_delay,
        addra_out     => FM_AAAA_L3PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L3PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L3PHIA_start
      );

    FM_BBBB_L3PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L3PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L3PHIA_wea_delay,
        addra     => FM_BBBB_L3PHIA_writeaddr_delay,
        dina      => FM_BBBB_L3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L3PHIA_V_readaddr,
        doutb     => FM_BBBB_L3PHIA_V_dout,
        sync_nent => FM_BBBB_L3PHIA_start,
        nent_o    => FM_BBBB_L3PHIA_AV_dout_nent
      );

    FM_BBBB_L3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L3PHIA_wea,
        addra     => FM_BBBB_L3PHIA_writeaddr,
        dina      => FM_BBBB_L3PHIA_din,
        wea_out       => FM_BBBB_L3PHIA_wea_delay,
        addra_out     => FM_BBBB_L3PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L3PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L3PHIA_start
      );

    FM_AAAA_L3PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L3PHIB_wea_delay,
        addra     => FM_AAAA_L3PHIB_writeaddr_delay,
        dina      => FM_AAAA_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L3PHIB_V_readaddr,
        doutb     => FM_AAAA_L3PHIB_V_dout,
        sync_nent => FM_AAAA_L3PHIB_start,
        nent_o    => FM_AAAA_L3PHIB_AV_dout_nent
      );

    FM_AAAA_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L3PHIB_wea,
        addra     => FM_AAAA_L3PHIB_writeaddr,
        dina      => FM_AAAA_L3PHIB_din,
        wea_out       => FM_AAAA_L3PHIB_wea_delay,
        addra_out     => FM_AAAA_L3PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L3PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L3PHIB_start
      );

    FM_BBBB_L3PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L3PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L3PHIB_wea_delay,
        addra     => FM_BBBB_L3PHIB_writeaddr_delay,
        dina      => FM_BBBB_L3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L3PHIB_V_readaddr,
        doutb     => FM_BBBB_L3PHIB_V_dout,
        sync_nent => FM_BBBB_L3PHIB_start,
        nent_o    => FM_BBBB_L3PHIB_AV_dout_nent
      );

    FM_BBBB_L3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L3PHIB_wea,
        addra     => FM_BBBB_L3PHIB_writeaddr,
        dina      => FM_BBBB_L3PHIB_din,
        wea_out       => FM_BBBB_L3PHIB_wea_delay,
        addra_out     => FM_BBBB_L3PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L3PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L3PHIB_start
      );

    FM_AAAA_L3PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L3PHIC_wea_delay,
        addra     => FM_AAAA_L3PHIC_writeaddr_delay,
        dina      => FM_AAAA_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L3PHIC_V_readaddr,
        doutb     => FM_AAAA_L3PHIC_V_dout,
        sync_nent => FM_AAAA_L3PHIC_start,
        nent_o    => FM_AAAA_L3PHIC_AV_dout_nent
      );

    FM_AAAA_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L3PHIC_wea,
        addra     => FM_AAAA_L3PHIC_writeaddr,
        dina      => FM_AAAA_L3PHIC_din,
        wea_out       => FM_AAAA_L3PHIC_wea_delay,
        addra_out     => FM_AAAA_L3PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L3PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L3PHIC_start
      );

    FM_BBBB_L3PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L3PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L3PHIC_wea_delay,
        addra     => FM_BBBB_L3PHIC_writeaddr_delay,
        dina      => FM_BBBB_L3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L3PHIC_V_readaddr,
        doutb     => FM_BBBB_L3PHIC_V_dout,
        sync_nent => FM_BBBB_L3PHIC_start,
        nent_o    => FM_BBBB_L3PHIC_AV_dout_nent
      );

    FM_BBBB_L3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L3PHIC_wea,
        addra     => FM_BBBB_L3PHIC_writeaddr,
        dina      => FM_BBBB_L3PHIC_din,
        wea_out       => FM_BBBB_L3PHIC_wea_delay,
        addra_out     => FM_BBBB_L3PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L3PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L3PHIC_start
      );

    FM_AAAA_L3PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L3PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L3PHID_wea_delay,
        addra     => FM_AAAA_L3PHID_writeaddr_delay,
        dina      => FM_AAAA_L3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L3PHID_V_readaddr,
        doutb     => FM_AAAA_L3PHID_V_dout,
        sync_nent => FM_AAAA_L3PHID_start,
        nent_o    => FM_AAAA_L3PHID_AV_dout_nent
      );

    FM_AAAA_L3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L3PHID_wea,
        addra     => FM_AAAA_L3PHID_writeaddr,
        dina      => FM_AAAA_L3PHID_din,
        wea_out       => FM_AAAA_L3PHID_wea_delay,
        addra_out     => FM_AAAA_L3PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L3PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L3PHID_start
      );

    FM_BBBB_L3PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L3PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L3PHID_wea_delay,
        addra     => FM_BBBB_L3PHID_writeaddr_delay,
        dina      => FM_BBBB_L3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L3PHID_V_readaddr,
        doutb     => FM_BBBB_L3PHID_V_dout,
        sync_nent => FM_BBBB_L3PHID_start,
        nent_o    => FM_BBBB_L3PHID_AV_dout_nent
      );

    FM_BBBB_L3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L3PHID_wea,
        addra     => FM_BBBB_L3PHID_writeaddr,
        dina      => FM_BBBB_L3PHID_din,
        wea_out       => FM_BBBB_L3PHID_wea_delay,
        addra_out     => FM_BBBB_L3PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L3PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L3PHID_start
      );

    FM_AAAA_L4PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L4PHIA_wea_delay,
        addra     => FM_AAAA_L4PHIA_writeaddr_delay,
        dina      => FM_AAAA_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L4PHIA_V_readaddr,
        doutb     => FM_AAAA_L4PHIA_V_dout,
        sync_nent => FM_AAAA_L4PHIA_start,
        nent_o    => FM_AAAA_L4PHIA_AV_dout_nent
      );

    FM_AAAA_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L4PHIA_wea,
        addra     => FM_AAAA_L4PHIA_writeaddr,
        dina      => FM_AAAA_L4PHIA_din,
        wea_out       => FM_AAAA_L4PHIA_wea_delay,
        addra_out     => FM_AAAA_L4PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L4PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L4PHIA_start
      );

    FM_BBBB_L4PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L4PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L4PHIA_wea_delay,
        addra     => FM_BBBB_L4PHIA_writeaddr_delay,
        dina      => FM_BBBB_L4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L4PHIA_V_readaddr,
        doutb     => FM_BBBB_L4PHIA_V_dout,
        sync_nent => FM_BBBB_L4PHIA_start,
        nent_o    => FM_BBBB_L4PHIA_AV_dout_nent
      );

    FM_BBBB_L4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L4PHIA_wea,
        addra     => FM_BBBB_L4PHIA_writeaddr,
        dina      => FM_BBBB_L4PHIA_din,
        wea_out       => FM_BBBB_L4PHIA_wea_delay,
        addra_out     => FM_BBBB_L4PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L4PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L4PHIA_start
      );

    FM_AAAA_L4PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L4PHIB_wea_delay,
        addra     => FM_AAAA_L4PHIB_writeaddr_delay,
        dina      => FM_AAAA_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L4PHIB_V_readaddr,
        doutb     => FM_AAAA_L4PHIB_V_dout,
        sync_nent => FM_AAAA_L4PHIB_start,
        nent_o    => FM_AAAA_L4PHIB_AV_dout_nent
      );

    FM_AAAA_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L4PHIB_wea,
        addra     => FM_AAAA_L4PHIB_writeaddr,
        dina      => FM_AAAA_L4PHIB_din,
        wea_out       => FM_AAAA_L4PHIB_wea_delay,
        addra_out     => FM_AAAA_L4PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L4PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L4PHIB_start
      );

    FM_BBBB_L4PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L4PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L4PHIB_wea_delay,
        addra     => FM_BBBB_L4PHIB_writeaddr_delay,
        dina      => FM_BBBB_L4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L4PHIB_V_readaddr,
        doutb     => FM_BBBB_L4PHIB_V_dout,
        sync_nent => FM_BBBB_L4PHIB_start,
        nent_o    => FM_BBBB_L4PHIB_AV_dout_nent
      );

    FM_BBBB_L4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L4PHIB_wea,
        addra     => FM_BBBB_L4PHIB_writeaddr,
        dina      => FM_BBBB_L4PHIB_din,
        wea_out       => FM_BBBB_L4PHIB_wea_delay,
        addra_out     => FM_BBBB_L4PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L4PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L4PHIB_start
      );

    FM_AAAA_L4PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L4PHIC_wea_delay,
        addra     => FM_AAAA_L4PHIC_writeaddr_delay,
        dina      => FM_AAAA_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L4PHIC_V_readaddr,
        doutb     => FM_AAAA_L4PHIC_V_dout,
        sync_nent => FM_AAAA_L4PHIC_start,
        nent_o    => FM_AAAA_L4PHIC_AV_dout_nent
      );

    FM_AAAA_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L4PHIC_wea,
        addra     => FM_AAAA_L4PHIC_writeaddr,
        dina      => FM_AAAA_L4PHIC_din,
        wea_out       => FM_AAAA_L4PHIC_wea_delay,
        addra_out     => FM_AAAA_L4PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L4PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L4PHIC_start
      );

    FM_BBBB_L4PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L4PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L4PHIC_wea_delay,
        addra     => FM_BBBB_L4PHIC_writeaddr_delay,
        dina      => FM_BBBB_L4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L4PHIC_V_readaddr,
        doutb     => FM_BBBB_L4PHIC_V_dout,
        sync_nent => FM_BBBB_L4PHIC_start,
        nent_o    => FM_BBBB_L4PHIC_AV_dout_nent
      );

    FM_BBBB_L4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L4PHIC_wea,
        addra     => FM_BBBB_L4PHIC_writeaddr,
        dina      => FM_BBBB_L4PHIC_din,
        wea_out       => FM_BBBB_L4PHIC_wea_delay,
        addra_out     => FM_BBBB_L4PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L4PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L4PHIC_start
      );

    FM_AAAA_L4PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L4PHID_wea_delay,
        addra     => FM_AAAA_L4PHID_writeaddr_delay,
        dina      => FM_AAAA_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L4PHID_V_readaddr,
        doutb     => FM_AAAA_L4PHID_V_dout,
        sync_nent => FM_AAAA_L4PHID_start,
        nent_o    => FM_AAAA_L4PHID_AV_dout_nent
      );

    FM_AAAA_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L4PHID_wea,
        addra     => FM_AAAA_L4PHID_writeaddr,
        dina      => FM_AAAA_L4PHID_din,
        wea_out       => FM_AAAA_L4PHID_wea_delay,
        addra_out     => FM_AAAA_L4PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L4PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L4PHID_start
      );

    FM_BBBB_L4PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L4PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L4PHID_wea_delay,
        addra     => FM_BBBB_L4PHID_writeaddr_delay,
        dina      => FM_BBBB_L4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L4PHID_V_readaddr,
        doutb     => FM_BBBB_L4PHID_V_dout,
        sync_nent => FM_BBBB_L4PHID_start,
        nent_o    => FM_BBBB_L4PHID_AV_dout_nent
      );

    FM_BBBB_L4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L4PHID_wea,
        addra     => FM_BBBB_L4PHID_writeaddr,
        dina      => FM_BBBB_L4PHID_din,
        wea_out       => FM_BBBB_L4PHID_wea_delay,
        addra_out     => FM_BBBB_L4PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L4PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L4PHID_start
      );

    FM_AAAA_L5PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L5PHIA_wea_delay,
        addra     => FM_AAAA_L5PHIA_writeaddr_delay,
        dina      => FM_AAAA_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L5PHIA_V_readaddr,
        doutb     => FM_AAAA_L5PHIA_V_dout,
        sync_nent => FM_AAAA_L5PHIA_start,
        nent_o    => FM_AAAA_L5PHIA_AV_dout_nent
      );

    FM_AAAA_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L5PHIA_wea,
        addra     => FM_AAAA_L5PHIA_writeaddr,
        dina      => FM_AAAA_L5PHIA_din,
        wea_out       => FM_AAAA_L5PHIA_wea_delay,
        addra_out     => FM_AAAA_L5PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L5PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L5PHIA_start
      );

    FM_BBBB_L5PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L5PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L5PHIA_wea_delay,
        addra     => FM_BBBB_L5PHIA_writeaddr_delay,
        dina      => FM_BBBB_L5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L5PHIA_V_readaddr,
        doutb     => FM_BBBB_L5PHIA_V_dout,
        sync_nent => FM_BBBB_L5PHIA_start,
        nent_o    => FM_BBBB_L5PHIA_AV_dout_nent
      );

    FM_BBBB_L5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L5PHIA_wea,
        addra     => FM_BBBB_L5PHIA_writeaddr,
        dina      => FM_BBBB_L5PHIA_din,
        wea_out       => FM_BBBB_L5PHIA_wea_delay,
        addra_out     => FM_BBBB_L5PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L5PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L5PHIA_start
      );

    FM_AAAA_L5PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L5PHIB_wea_delay,
        addra     => FM_AAAA_L5PHIB_writeaddr_delay,
        dina      => FM_AAAA_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L5PHIB_V_readaddr,
        doutb     => FM_AAAA_L5PHIB_V_dout,
        sync_nent => FM_AAAA_L5PHIB_start,
        nent_o    => FM_AAAA_L5PHIB_AV_dout_nent
      );

    FM_AAAA_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L5PHIB_wea,
        addra     => FM_AAAA_L5PHIB_writeaddr,
        dina      => FM_AAAA_L5PHIB_din,
        wea_out       => FM_AAAA_L5PHIB_wea_delay,
        addra_out     => FM_AAAA_L5PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L5PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L5PHIB_start
      );

    FM_BBBB_L5PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L5PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L5PHIB_wea_delay,
        addra     => FM_BBBB_L5PHIB_writeaddr_delay,
        dina      => FM_BBBB_L5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L5PHIB_V_readaddr,
        doutb     => FM_BBBB_L5PHIB_V_dout,
        sync_nent => FM_BBBB_L5PHIB_start,
        nent_o    => FM_BBBB_L5PHIB_AV_dout_nent
      );

    FM_BBBB_L5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L5PHIB_wea,
        addra     => FM_BBBB_L5PHIB_writeaddr,
        dina      => FM_BBBB_L5PHIB_din,
        wea_out       => FM_BBBB_L5PHIB_wea_delay,
        addra_out     => FM_BBBB_L5PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L5PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L5PHIB_start
      );

    FM_AAAA_L5PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L5PHIC_wea_delay,
        addra     => FM_AAAA_L5PHIC_writeaddr_delay,
        dina      => FM_AAAA_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L5PHIC_V_readaddr,
        doutb     => FM_AAAA_L5PHIC_V_dout,
        sync_nent => FM_AAAA_L5PHIC_start,
        nent_o    => FM_AAAA_L5PHIC_AV_dout_nent
      );

    FM_AAAA_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L5PHIC_wea,
        addra     => FM_AAAA_L5PHIC_writeaddr,
        dina      => FM_AAAA_L5PHIC_din,
        wea_out       => FM_AAAA_L5PHIC_wea_delay,
        addra_out     => FM_AAAA_L5PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L5PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L5PHIC_start
      );

    FM_BBBB_L5PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L5PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L5PHIC_wea_delay,
        addra     => FM_BBBB_L5PHIC_writeaddr_delay,
        dina      => FM_BBBB_L5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L5PHIC_V_readaddr,
        doutb     => FM_BBBB_L5PHIC_V_dout,
        sync_nent => FM_BBBB_L5PHIC_start,
        nent_o    => FM_BBBB_L5PHIC_AV_dout_nent
      );

    FM_BBBB_L5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L5PHIC_wea,
        addra     => FM_BBBB_L5PHIC_writeaddr,
        dina      => FM_BBBB_L5PHIC_din,
        wea_out       => FM_BBBB_L5PHIC_wea_delay,
        addra_out     => FM_BBBB_L5PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L5PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L5PHIC_start
      );

    FM_AAAA_L5PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L5PHID_wea_delay,
        addra     => FM_AAAA_L5PHID_writeaddr_delay,
        dina      => FM_AAAA_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L5PHID_V_readaddr,
        doutb     => FM_AAAA_L5PHID_V_dout,
        sync_nent => FM_AAAA_L5PHID_start,
        nent_o    => FM_AAAA_L5PHID_AV_dout_nent
      );

    FM_AAAA_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L5PHID_wea,
        addra     => FM_AAAA_L5PHID_writeaddr,
        dina      => FM_AAAA_L5PHID_din,
        wea_out       => FM_AAAA_L5PHID_wea_delay,
        addra_out     => FM_AAAA_L5PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L5PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L5PHID_start
      );

    FM_BBBB_L5PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L5PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L5PHID_wea_delay,
        addra     => FM_BBBB_L5PHID_writeaddr_delay,
        dina      => FM_BBBB_L5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L5PHID_V_readaddr,
        doutb     => FM_BBBB_L5PHID_V_dout,
        sync_nent => FM_BBBB_L5PHID_start,
        nent_o    => FM_BBBB_L5PHID_AV_dout_nent
      );

    FM_BBBB_L5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L5PHID_wea,
        addra     => FM_BBBB_L5PHID_writeaddr,
        dina      => FM_BBBB_L5PHID_din,
        wea_out       => FM_BBBB_L5PHID_wea_delay,
        addra_out     => FM_BBBB_L5PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L5PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L5PHID_start
      );

    FM_AAAA_L6PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L6PHIA_wea_delay,
        addra     => FM_AAAA_L6PHIA_writeaddr_delay,
        dina      => FM_AAAA_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L6PHIA_V_readaddr,
        doutb     => FM_AAAA_L6PHIA_V_dout,
        sync_nent => FM_AAAA_L6PHIA_start,
        nent_o    => FM_AAAA_L6PHIA_AV_dout_nent
      );

    FM_AAAA_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L6PHIA_wea,
        addra     => FM_AAAA_L6PHIA_writeaddr,
        dina      => FM_AAAA_L6PHIA_din,
        wea_out       => FM_AAAA_L6PHIA_wea_delay,
        addra_out     => FM_AAAA_L6PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_L6PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L6PHIA_start
      );

    FM_BBBB_L6PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L6PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L6PHIA_wea_delay,
        addra     => FM_BBBB_L6PHIA_writeaddr_delay,
        dina      => FM_BBBB_L6PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L6PHIA_V_readaddr,
        doutb     => FM_BBBB_L6PHIA_V_dout,
        sync_nent => FM_BBBB_L6PHIA_start,
        nent_o    => FM_BBBB_L6PHIA_AV_dout_nent
      );

    FM_BBBB_L6PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L6PHIA_wea,
        addra     => FM_BBBB_L6PHIA_writeaddr,
        dina      => FM_BBBB_L6PHIA_din,
        wea_out       => FM_BBBB_L6PHIA_wea_delay,
        addra_out     => FM_BBBB_L6PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_L6PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L6PHIA_start
      );

    FM_AAAA_L6PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L6PHIB_wea_delay,
        addra     => FM_AAAA_L6PHIB_writeaddr_delay,
        dina      => FM_AAAA_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L6PHIB_V_readaddr,
        doutb     => FM_AAAA_L6PHIB_V_dout,
        sync_nent => FM_AAAA_L6PHIB_start,
        nent_o    => FM_AAAA_L6PHIB_AV_dout_nent
      );

    FM_AAAA_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L6PHIB_wea,
        addra     => FM_AAAA_L6PHIB_writeaddr,
        dina      => FM_AAAA_L6PHIB_din,
        wea_out       => FM_AAAA_L6PHIB_wea_delay,
        addra_out     => FM_AAAA_L6PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_L6PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L6PHIB_start
      );

    FM_BBBB_L6PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L6PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L6PHIB_wea_delay,
        addra     => FM_BBBB_L6PHIB_writeaddr_delay,
        dina      => FM_BBBB_L6PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L6PHIB_V_readaddr,
        doutb     => FM_BBBB_L6PHIB_V_dout,
        sync_nent => FM_BBBB_L6PHIB_start,
        nent_o    => FM_BBBB_L6PHIB_AV_dout_nent
      );

    FM_BBBB_L6PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L6PHIB_wea,
        addra     => FM_BBBB_L6PHIB_writeaddr,
        dina      => FM_BBBB_L6PHIB_din,
        wea_out       => FM_BBBB_L6PHIB_wea_delay,
        addra_out     => FM_BBBB_L6PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_L6PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L6PHIB_start
      );

    FM_AAAA_L6PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L6PHIC_wea_delay,
        addra     => FM_AAAA_L6PHIC_writeaddr_delay,
        dina      => FM_AAAA_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L6PHIC_V_readaddr,
        doutb     => FM_AAAA_L6PHIC_V_dout,
        sync_nent => FM_AAAA_L6PHIC_start,
        nent_o    => FM_AAAA_L6PHIC_AV_dout_nent
      );

    FM_AAAA_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L6PHIC_wea,
        addra     => FM_AAAA_L6PHIC_writeaddr,
        dina      => FM_AAAA_L6PHIC_din,
        wea_out       => FM_AAAA_L6PHIC_wea_delay,
        addra_out     => FM_AAAA_L6PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_L6PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L6PHIC_start
      );

    FM_BBBB_L6PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L6PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L6PHIC_wea_delay,
        addra     => FM_BBBB_L6PHIC_writeaddr_delay,
        dina      => FM_BBBB_L6PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L6PHIC_V_readaddr,
        doutb     => FM_BBBB_L6PHIC_V_dout,
        sync_nent => FM_BBBB_L6PHIC_start,
        nent_o    => FM_BBBB_L6PHIC_AV_dout_nent
      );

    FM_BBBB_L6PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L6PHIC_wea,
        addra     => FM_BBBB_L6PHIC_writeaddr,
        dina      => FM_BBBB_L6PHIC_din,
        wea_out       => FM_BBBB_L6PHIC_wea_delay,
        addra_out     => FM_BBBB_L6PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_L6PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L6PHIC_start
      );

    FM_AAAA_L6PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_L6PHID_wea_delay,
        addra     => FM_AAAA_L6PHID_writeaddr_delay,
        dina      => FM_AAAA_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_L6PHID_V_readaddr,
        doutb     => FM_AAAA_L6PHID_V_dout,
        sync_nent => FM_AAAA_L6PHID_start,
        nent_o    => FM_AAAA_L6PHID_AV_dout_nent
      );

    FM_AAAA_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_L6PHID_wea,
        addra     => FM_AAAA_L6PHID_writeaddr,
        dina      => FM_AAAA_L6PHID_din,
        wea_out       => FM_AAAA_L6PHID_wea_delay,
        addra_out     => FM_AAAA_L6PHID_writeaddr_delay,
        dina_out      => FM_AAAA_L6PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_L6PHID_start
      );

    FM_BBBB_L6PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 52,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_L6PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_L6PHID_wea_delay,
        addra     => FM_BBBB_L6PHID_writeaddr_delay,
        dina      => FM_BBBB_L6PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_L6PHID_V_readaddr,
        doutb     => FM_BBBB_L6PHID_V_dout,
        sync_nent => FM_BBBB_L6PHID_start,
        nent_o    => FM_BBBB_L6PHID_AV_dout_nent
      );

    FM_BBBB_L6PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 52
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_L6PHID_wea,
        addra     => FM_BBBB_L6PHID_writeaddr,
        dina      => FM_BBBB_L6PHID_din,
        wea_out       => FM_BBBB_L6PHID_wea_delay,
        addra_out     => FM_BBBB_L6PHID_writeaddr_delay,
        dina_out      => FM_BBBB_L6PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_L6PHID_start
      );

    FM_AAAA_D1PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D1PHIA_wea_delay,
        addra     => FM_AAAA_D1PHIA_writeaddr_delay,
        dina      => FM_AAAA_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D1PHIA_V_readaddr,
        doutb     => FM_AAAA_D1PHIA_V_dout,
        sync_nent => FM_AAAA_D1PHIA_start,
        nent_o    => FM_AAAA_D1PHIA_AV_dout_nent
      );

    FM_AAAA_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D1PHIA_wea,
        addra     => FM_AAAA_D1PHIA_writeaddr,
        dina      => FM_AAAA_D1PHIA_din,
        wea_out       => FM_AAAA_D1PHIA_wea_delay,
        addra_out     => FM_AAAA_D1PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_D1PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D1PHIA_start
      );

    FM_BBBB_D1PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D1PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D1PHIA_wea_delay,
        addra     => FM_BBBB_D1PHIA_writeaddr_delay,
        dina      => FM_BBBB_D1PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D1PHIA_V_readaddr,
        doutb     => FM_BBBB_D1PHIA_V_dout,
        sync_nent => FM_BBBB_D1PHIA_start,
        nent_o    => FM_BBBB_D1PHIA_AV_dout_nent
      );

    FM_BBBB_D1PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D1PHIA_wea,
        addra     => FM_BBBB_D1PHIA_writeaddr,
        dina      => FM_BBBB_D1PHIA_din,
        wea_out       => FM_BBBB_D1PHIA_wea_delay,
        addra_out     => FM_BBBB_D1PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_D1PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D1PHIA_start
      );

    FM_AAAA_D1PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D1PHIB_wea_delay,
        addra     => FM_AAAA_D1PHIB_writeaddr_delay,
        dina      => FM_AAAA_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D1PHIB_V_readaddr,
        doutb     => FM_AAAA_D1PHIB_V_dout,
        sync_nent => FM_AAAA_D1PHIB_start,
        nent_o    => FM_AAAA_D1PHIB_AV_dout_nent
      );

    FM_AAAA_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D1PHIB_wea,
        addra     => FM_AAAA_D1PHIB_writeaddr,
        dina      => FM_AAAA_D1PHIB_din,
        wea_out       => FM_AAAA_D1PHIB_wea_delay,
        addra_out     => FM_AAAA_D1PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_D1PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D1PHIB_start
      );

    FM_BBBB_D1PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D1PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D1PHIB_wea_delay,
        addra     => FM_BBBB_D1PHIB_writeaddr_delay,
        dina      => FM_BBBB_D1PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D1PHIB_V_readaddr,
        doutb     => FM_BBBB_D1PHIB_V_dout,
        sync_nent => FM_BBBB_D1PHIB_start,
        nent_o    => FM_BBBB_D1PHIB_AV_dout_nent
      );

    FM_BBBB_D1PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D1PHIB_wea,
        addra     => FM_BBBB_D1PHIB_writeaddr,
        dina      => FM_BBBB_D1PHIB_din,
        wea_out       => FM_BBBB_D1PHIB_wea_delay,
        addra_out     => FM_BBBB_D1PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_D1PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D1PHIB_start
      );

    FM_AAAA_D1PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D1PHIC_wea_delay,
        addra     => FM_AAAA_D1PHIC_writeaddr_delay,
        dina      => FM_AAAA_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D1PHIC_V_readaddr,
        doutb     => FM_AAAA_D1PHIC_V_dout,
        sync_nent => FM_AAAA_D1PHIC_start,
        nent_o    => FM_AAAA_D1PHIC_AV_dout_nent
      );

    FM_AAAA_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D1PHIC_wea,
        addra     => FM_AAAA_D1PHIC_writeaddr,
        dina      => FM_AAAA_D1PHIC_din,
        wea_out       => FM_AAAA_D1PHIC_wea_delay,
        addra_out     => FM_AAAA_D1PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_D1PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D1PHIC_start
      );

    FM_BBBB_D1PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D1PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D1PHIC_wea_delay,
        addra     => FM_BBBB_D1PHIC_writeaddr_delay,
        dina      => FM_BBBB_D1PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D1PHIC_V_readaddr,
        doutb     => FM_BBBB_D1PHIC_V_dout,
        sync_nent => FM_BBBB_D1PHIC_start,
        nent_o    => FM_BBBB_D1PHIC_AV_dout_nent
      );

    FM_BBBB_D1PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D1PHIC_wea,
        addra     => FM_BBBB_D1PHIC_writeaddr,
        dina      => FM_BBBB_D1PHIC_din,
        wea_out       => FM_BBBB_D1PHIC_wea_delay,
        addra_out     => FM_BBBB_D1PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_D1PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D1PHIC_start
      );

    FM_AAAA_D1PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D1PHID_wea_delay,
        addra     => FM_AAAA_D1PHID_writeaddr_delay,
        dina      => FM_AAAA_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D1PHID_V_readaddr,
        doutb     => FM_AAAA_D1PHID_V_dout,
        sync_nent => FM_AAAA_D1PHID_start,
        nent_o    => FM_AAAA_D1PHID_AV_dout_nent
      );

    FM_AAAA_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D1PHID_wea,
        addra     => FM_AAAA_D1PHID_writeaddr,
        dina      => FM_AAAA_D1PHID_din,
        wea_out       => FM_AAAA_D1PHID_wea_delay,
        addra_out     => FM_AAAA_D1PHID_writeaddr_delay,
        dina_out      => FM_AAAA_D1PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D1PHID_start
      );

    FM_BBBB_D1PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D1PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D1PHID_wea_delay,
        addra     => FM_BBBB_D1PHID_writeaddr_delay,
        dina      => FM_BBBB_D1PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D1PHID_V_readaddr,
        doutb     => FM_BBBB_D1PHID_V_dout,
        sync_nent => FM_BBBB_D1PHID_start,
        nent_o    => FM_BBBB_D1PHID_AV_dout_nent
      );

    FM_BBBB_D1PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D1PHID_wea,
        addra     => FM_BBBB_D1PHID_writeaddr,
        dina      => FM_BBBB_D1PHID_din,
        wea_out       => FM_BBBB_D1PHID_wea_delay,
        addra_out     => FM_BBBB_D1PHID_writeaddr_delay,
        dina_out      => FM_BBBB_D1PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D1PHID_start
      );

    FM_AAAA_D2PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D2PHIA_wea_delay,
        addra     => FM_AAAA_D2PHIA_writeaddr_delay,
        dina      => FM_AAAA_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D2PHIA_V_readaddr,
        doutb     => FM_AAAA_D2PHIA_V_dout,
        sync_nent => FM_AAAA_D2PHIA_start,
        nent_o    => FM_AAAA_D2PHIA_AV_dout_nent
      );

    FM_AAAA_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D2PHIA_wea,
        addra     => FM_AAAA_D2PHIA_writeaddr,
        dina      => FM_AAAA_D2PHIA_din,
        wea_out       => FM_AAAA_D2PHIA_wea_delay,
        addra_out     => FM_AAAA_D2PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_D2PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D2PHIA_start
      );

    FM_BBBB_D2PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D2PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D2PHIA_wea_delay,
        addra     => FM_BBBB_D2PHIA_writeaddr_delay,
        dina      => FM_BBBB_D2PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D2PHIA_V_readaddr,
        doutb     => FM_BBBB_D2PHIA_V_dout,
        sync_nent => FM_BBBB_D2PHIA_start,
        nent_o    => FM_BBBB_D2PHIA_AV_dout_nent
      );

    FM_BBBB_D2PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D2PHIA_wea,
        addra     => FM_BBBB_D2PHIA_writeaddr,
        dina      => FM_BBBB_D2PHIA_din,
        wea_out       => FM_BBBB_D2PHIA_wea_delay,
        addra_out     => FM_BBBB_D2PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_D2PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D2PHIA_start
      );

    FM_AAAA_D2PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D2PHIB_wea_delay,
        addra     => FM_AAAA_D2PHIB_writeaddr_delay,
        dina      => FM_AAAA_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D2PHIB_V_readaddr,
        doutb     => FM_AAAA_D2PHIB_V_dout,
        sync_nent => FM_AAAA_D2PHIB_start,
        nent_o    => FM_AAAA_D2PHIB_AV_dout_nent
      );

    FM_AAAA_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D2PHIB_wea,
        addra     => FM_AAAA_D2PHIB_writeaddr,
        dina      => FM_AAAA_D2PHIB_din,
        wea_out       => FM_AAAA_D2PHIB_wea_delay,
        addra_out     => FM_AAAA_D2PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_D2PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D2PHIB_start
      );

    FM_BBBB_D2PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D2PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D2PHIB_wea_delay,
        addra     => FM_BBBB_D2PHIB_writeaddr_delay,
        dina      => FM_BBBB_D2PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D2PHIB_V_readaddr,
        doutb     => FM_BBBB_D2PHIB_V_dout,
        sync_nent => FM_BBBB_D2PHIB_start,
        nent_o    => FM_BBBB_D2PHIB_AV_dout_nent
      );

    FM_BBBB_D2PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D2PHIB_wea,
        addra     => FM_BBBB_D2PHIB_writeaddr,
        dina      => FM_BBBB_D2PHIB_din,
        wea_out       => FM_BBBB_D2PHIB_wea_delay,
        addra_out     => FM_BBBB_D2PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_D2PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D2PHIB_start
      );

    FM_AAAA_D2PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D2PHIC_wea_delay,
        addra     => FM_AAAA_D2PHIC_writeaddr_delay,
        dina      => FM_AAAA_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D2PHIC_V_readaddr,
        doutb     => FM_AAAA_D2PHIC_V_dout,
        sync_nent => FM_AAAA_D2PHIC_start,
        nent_o    => FM_AAAA_D2PHIC_AV_dout_nent
      );

    FM_AAAA_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D2PHIC_wea,
        addra     => FM_AAAA_D2PHIC_writeaddr,
        dina      => FM_AAAA_D2PHIC_din,
        wea_out       => FM_AAAA_D2PHIC_wea_delay,
        addra_out     => FM_AAAA_D2PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_D2PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D2PHIC_start
      );

    FM_BBBB_D2PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D2PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D2PHIC_wea_delay,
        addra     => FM_BBBB_D2PHIC_writeaddr_delay,
        dina      => FM_BBBB_D2PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D2PHIC_V_readaddr,
        doutb     => FM_BBBB_D2PHIC_V_dout,
        sync_nent => FM_BBBB_D2PHIC_start,
        nent_o    => FM_BBBB_D2PHIC_AV_dout_nent
      );

    FM_BBBB_D2PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D2PHIC_wea,
        addra     => FM_BBBB_D2PHIC_writeaddr,
        dina      => FM_BBBB_D2PHIC_din,
        wea_out       => FM_BBBB_D2PHIC_wea_delay,
        addra_out     => FM_BBBB_D2PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_D2PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D2PHIC_start
      );

    FM_AAAA_D2PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D2PHID_wea_delay,
        addra     => FM_AAAA_D2PHID_writeaddr_delay,
        dina      => FM_AAAA_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D2PHID_V_readaddr,
        doutb     => FM_AAAA_D2PHID_V_dout,
        sync_nent => FM_AAAA_D2PHID_start,
        nent_o    => FM_AAAA_D2PHID_AV_dout_nent
      );

    FM_AAAA_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D2PHID_wea,
        addra     => FM_AAAA_D2PHID_writeaddr,
        dina      => FM_AAAA_D2PHID_din,
        wea_out       => FM_AAAA_D2PHID_wea_delay,
        addra_out     => FM_AAAA_D2PHID_writeaddr_delay,
        dina_out      => FM_AAAA_D2PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D2PHID_start
      );

    FM_BBBB_D2PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D2PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D2PHID_wea_delay,
        addra     => FM_BBBB_D2PHID_writeaddr_delay,
        dina      => FM_BBBB_D2PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D2PHID_V_readaddr,
        doutb     => FM_BBBB_D2PHID_V_dout,
        sync_nent => FM_BBBB_D2PHID_start,
        nent_o    => FM_BBBB_D2PHID_AV_dout_nent
      );

    FM_BBBB_D2PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D2PHID_wea,
        addra     => FM_BBBB_D2PHID_writeaddr,
        dina      => FM_BBBB_D2PHID_din,
        wea_out       => FM_BBBB_D2PHID_wea_delay,
        addra_out     => FM_BBBB_D2PHID_writeaddr_delay,
        dina_out      => FM_BBBB_D2PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D2PHID_start
      );

    FM_AAAA_D3PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D3PHIA_wea_delay,
        addra     => FM_AAAA_D3PHIA_writeaddr_delay,
        dina      => FM_AAAA_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D3PHIA_V_readaddr,
        doutb     => FM_AAAA_D3PHIA_V_dout,
        sync_nent => FM_AAAA_D3PHIA_start,
        nent_o    => FM_AAAA_D3PHIA_AV_dout_nent
      );

    FM_AAAA_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D3PHIA_wea,
        addra     => FM_AAAA_D3PHIA_writeaddr,
        dina      => FM_AAAA_D3PHIA_din,
        wea_out       => FM_AAAA_D3PHIA_wea_delay,
        addra_out     => FM_AAAA_D3PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_D3PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D3PHIA_start
      );

    FM_BBBB_D3PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D3PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D3PHIA_wea_delay,
        addra     => FM_BBBB_D3PHIA_writeaddr_delay,
        dina      => FM_BBBB_D3PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D3PHIA_V_readaddr,
        doutb     => FM_BBBB_D3PHIA_V_dout,
        sync_nent => FM_BBBB_D3PHIA_start,
        nent_o    => FM_BBBB_D3PHIA_AV_dout_nent
      );

    FM_BBBB_D3PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D3PHIA_wea,
        addra     => FM_BBBB_D3PHIA_writeaddr,
        dina      => FM_BBBB_D3PHIA_din,
        wea_out       => FM_BBBB_D3PHIA_wea_delay,
        addra_out     => FM_BBBB_D3PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_D3PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D3PHIA_start
      );

    FM_AAAA_D3PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D3PHIB_wea_delay,
        addra     => FM_AAAA_D3PHIB_writeaddr_delay,
        dina      => FM_AAAA_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D3PHIB_V_readaddr,
        doutb     => FM_AAAA_D3PHIB_V_dout,
        sync_nent => FM_AAAA_D3PHIB_start,
        nent_o    => FM_AAAA_D3PHIB_AV_dout_nent
      );

    FM_AAAA_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D3PHIB_wea,
        addra     => FM_AAAA_D3PHIB_writeaddr,
        dina      => FM_AAAA_D3PHIB_din,
        wea_out       => FM_AAAA_D3PHIB_wea_delay,
        addra_out     => FM_AAAA_D3PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_D3PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D3PHIB_start
      );

    FM_BBBB_D3PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D3PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D3PHIB_wea_delay,
        addra     => FM_BBBB_D3PHIB_writeaddr_delay,
        dina      => FM_BBBB_D3PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D3PHIB_V_readaddr,
        doutb     => FM_BBBB_D3PHIB_V_dout,
        sync_nent => FM_BBBB_D3PHIB_start,
        nent_o    => FM_BBBB_D3PHIB_AV_dout_nent
      );

    FM_BBBB_D3PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D3PHIB_wea,
        addra     => FM_BBBB_D3PHIB_writeaddr,
        dina      => FM_BBBB_D3PHIB_din,
        wea_out       => FM_BBBB_D3PHIB_wea_delay,
        addra_out     => FM_BBBB_D3PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_D3PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D3PHIB_start
      );

    FM_AAAA_D3PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D3PHIC_wea_delay,
        addra     => FM_AAAA_D3PHIC_writeaddr_delay,
        dina      => FM_AAAA_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D3PHIC_V_readaddr,
        doutb     => FM_AAAA_D3PHIC_V_dout,
        sync_nent => FM_AAAA_D3PHIC_start,
        nent_o    => FM_AAAA_D3PHIC_AV_dout_nent
      );

    FM_AAAA_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D3PHIC_wea,
        addra     => FM_AAAA_D3PHIC_writeaddr,
        dina      => FM_AAAA_D3PHIC_din,
        wea_out       => FM_AAAA_D3PHIC_wea_delay,
        addra_out     => FM_AAAA_D3PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_D3PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D3PHIC_start
      );

    FM_BBBB_D3PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D3PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D3PHIC_wea_delay,
        addra     => FM_BBBB_D3PHIC_writeaddr_delay,
        dina      => FM_BBBB_D3PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D3PHIC_V_readaddr,
        doutb     => FM_BBBB_D3PHIC_V_dout,
        sync_nent => FM_BBBB_D3PHIC_start,
        nent_o    => FM_BBBB_D3PHIC_AV_dout_nent
      );

    FM_BBBB_D3PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D3PHIC_wea,
        addra     => FM_BBBB_D3PHIC_writeaddr,
        dina      => FM_BBBB_D3PHIC_din,
        wea_out       => FM_BBBB_D3PHIC_wea_delay,
        addra_out     => FM_BBBB_D3PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_D3PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D3PHIC_start
      );

    FM_AAAA_D3PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D3PHID_wea_delay,
        addra     => FM_AAAA_D3PHID_writeaddr_delay,
        dina      => FM_AAAA_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D3PHID_V_readaddr,
        doutb     => FM_AAAA_D3PHID_V_dout,
        sync_nent => FM_AAAA_D3PHID_start,
        nent_o    => FM_AAAA_D3PHID_AV_dout_nent
      );

    FM_AAAA_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D3PHID_wea,
        addra     => FM_AAAA_D3PHID_writeaddr,
        dina      => FM_AAAA_D3PHID_din,
        wea_out       => FM_AAAA_D3PHID_wea_delay,
        addra_out     => FM_AAAA_D3PHID_writeaddr_delay,
        dina_out      => FM_AAAA_D3PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D3PHID_start
      );

    FM_BBBB_D3PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D3PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D3PHID_wea_delay,
        addra     => FM_BBBB_D3PHID_writeaddr_delay,
        dina      => FM_BBBB_D3PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D3PHID_V_readaddr,
        doutb     => FM_BBBB_D3PHID_V_dout,
        sync_nent => FM_BBBB_D3PHID_start,
        nent_o    => FM_BBBB_D3PHID_AV_dout_nent
      );

    FM_BBBB_D3PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D3PHID_wea,
        addra     => FM_BBBB_D3PHID_writeaddr,
        dina      => FM_BBBB_D3PHID_din,
        wea_out       => FM_BBBB_D3PHID_wea_delay,
        addra_out     => FM_BBBB_D3PHID_writeaddr_delay,
        dina_out      => FM_BBBB_D3PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D3PHID_start
      );

    FM_AAAA_D4PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D4PHIA_wea_delay,
        addra     => FM_AAAA_D4PHIA_writeaddr_delay,
        dina      => FM_AAAA_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D4PHIA_V_readaddr,
        doutb     => FM_AAAA_D4PHIA_V_dout,
        sync_nent => FM_AAAA_D4PHIA_start,
        nent_o    => FM_AAAA_D4PHIA_AV_dout_nent
      );

    FM_AAAA_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D4PHIA_wea,
        addra     => FM_AAAA_D4PHIA_writeaddr,
        dina      => FM_AAAA_D4PHIA_din,
        wea_out       => FM_AAAA_D4PHIA_wea_delay,
        addra_out     => FM_AAAA_D4PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_D4PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D4PHIA_start
      );

    FM_BBBB_D4PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D4PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D4PHIA_wea_delay,
        addra     => FM_BBBB_D4PHIA_writeaddr_delay,
        dina      => FM_BBBB_D4PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D4PHIA_V_readaddr,
        doutb     => FM_BBBB_D4PHIA_V_dout,
        sync_nent => FM_BBBB_D4PHIA_start,
        nent_o    => FM_BBBB_D4PHIA_AV_dout_nent
      );

    FM_BBBB_D4PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D4PHIA_wea,
        addra     => FM_BBBB_D4PHIA_writeaddr,
        dina      => FM_BBBB_D4PHIA_din,
        wea_out       => FM_BBBB_D4PHIA_wea_delay,
        addra_out     => FM_BBBB_D4PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_D4PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D4PHIA_start
      );

    FM_AAAA_D4PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D4PHIB_wea_delay,
        addra     => FM_AAAA_D4PHIB_writeaddr_delay,
        dina      => FM_AAAA_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D4PHIB_V_readaddr,
        doutb     => FM_AAAA_D4PHIB_V_dout,
        sync_nent => FM_AAAA_D4PHIB_start,
        nent_o    => FM_AAAA_D4PHIB_AV_dout_nent
      );

    FM_AAAA_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D4PHIB_wea,
        addra     => FM_AAAA_D4PHIB_writeaddr,
        dina      => FM_AAAA_D4PHIB_din,
        wea_out       => FM_AAAA_D4PHIB_wea_delay,
        addra_out     => FM_AAAA_D4PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_D4PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D4PHIB_start
      );

    FM_BBBB_D4PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D4PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D4PHIB_wea_delay,
        addra     => FM_BBBB_D4PHIB_writeaddr_delay,
        dina      => FM_BBBB_D4PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D4PHIB_V_readaddr,
        doutb     => FM_BBBB_D4PHIB_V_dout,
        sync_nent => FM_BBBB_D4PHIB_start,
        nent_o    => FM_BBBB_D4PHIB_AV_dout_nent
      );

    FM_BBBB_D4PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D4PHIB_wea,
        addra     => FM_BBBB_D4PHIB_writeaddr,
        dina      => FM_BBBB_D4PHIB_din,
        wea_out       => FM_BBBB_D4PHIB_wea_delay,
        addra_out     => FM_BBBB_D4PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_D4PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D4PHIB_start
      );

    FM_AAAA_D4PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D4PHIC_wea_delay,
        addra     => FM_AAAA_D4PHIC_writeaddr_delay,
        dina      => FM_AAAA_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D4PHIC_V_readaddr,
        doutb     => FM_AAAA_D4PHIC_V_dout,
        sync_nent => FM_AAAA_D4PHIC_start,
        nent_o    => FM_AAAA_D4PHIC_AV_dout_nent
      );

    FM_AAAA_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D4PHIC_wea,
        addra     => FM_AAAA_D4PHIC_writeaddr,
        dina      => FM_AAAA_D4PHIC_din,
        wea_out       => FM_AAAA_D4PHIC_wea_delay,
        addra_out     => FM_AAAA_D4PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_D4PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D4PHIC_start
      );

    FM_BBBB_D4PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D4PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D4PHIC_wea_delay,
        addra     => FM_BBBB_D4PHIC_writeaddr_delay,
        dina      => FM_BBBB_D4PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D4PHIC_V_readaddr,
        doutb     => FM_BBBB_D4PHIC_V_dout,
        sync_nent => FM_BBBB_D4PHIC_start,
        nent_o    => FM_BBBB_D4PHIC_AV_dout_nent
      );

    FM_BBBB_D4PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D4PHIC_wea,
        addra     => FM_BBBB_D4PHIC_writeaddr,
        dina      => FM_BBBB_D4PHIC_din,
        wea_out       => FM_BBBB_D4PHIC_wea_delay,
        addra_out     => FM_BBBB_D4PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_D4PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D4PHIC_start
      );

    FM_AAAA_D4PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D4PHID_wea_delay,
        addra     => FM_AAAA_D4PHID_writeaddr_delay,
        dina      => FM_AAAA_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D4PHID_V_readaddr,
        doutb     => FM_AAAA_D4PHID_V_dout,
        sync_nent => FM_AAAA_D4PHID_start,
        nent_o    => FM_AAAA_D4PHID_AV_dout_nent
      );

    FM_AAAA_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D4PHID_wea,
        addra     => FM_AAAA_D4PHID_writeaddr,
        dina      => FM_AAAA_D4PHID_din,
        wea_out       => FM_AAAA_D4PHID_wea_delay,
        addra_out     => FM_AAAA_D4PHID_writeaddr_delay,
        dina_out      => FM_AAAA_D4PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D4PHID_start
      );

    FM_BBBB_D4PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D4PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D4PHID_wea_delay,
        addra     => FM_BBBB_D4PHID_writeaddr_delay,
        dina      => FM_BBBB_D4PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D4PHID_V_readaddr,
        doutb     => FM_BBBB_D4PHID_V_dout,
        sync_nent => FM_BBBB_D4PHID_start,
        nent_o    => FM_BBBB_D4PHID_AV_dout_nent
      );

    FM_BBBB_D4PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D4PHID_wea,
        addra     => FM_BBBB_D4PHID_writeaddr,
        dina      => FM_BBBB_D4PHID_din,
        wea_out       => FM_BBBB_D4PHID_wea_delay,
        addra_out     => FM_BBBB_D4PHID_writeaddr_delay,
        dina_out      => FM_BBBB_D4PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D4PHID_start
      );

    FM_AAAA_D5PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D5PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D5PHIA_wea_delay,
        addra     => FM_AAAA_D5PHIA_writeaddr_delay,
        dina      => FM_AAAA_D5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D5PHIA_V_readaddr,
        doutb     => FM_AAAA_D5PHIA_V_dout,
        sync_nent => FM_AAAA_D5PHIA_start,
        nent_o    => FM_AAAA_D5PHIA_AV_dout_nent
      );

    FM_AAAA_D5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D5PHIA_wea,
        addra     => FM_AAAA_D5PHIA_writeaddr,
        dina      => FM_AAAA_D5PHIA_din,
        wea_out       => FM_AAAA_D5PHIA_wea_delay,
        addra_out     => FM_AAAA_D5PHIA_writeaddr_delay,
        dina_out      => FM_AAAA_D5PHIA_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D5PHIA_start
      );

    FM_BBBB_D5PHIA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D5PHIA"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D5PHIA_wea_delay,
        addra     => FM_BBBB_D5PHIA_writeaddr_delay,
        dina      => FM_BBBB_D5PHIA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D5PHIA_V_readaddr,
        doutb     => FM_BBBB_D5PHIA_V_dout,
        sync_nent => FM_BBBB_D5PHIA_start,
        nent_o    => FM_BBBB_D5PHIA_AV_dout_nent
      );

    FM_BBBB_D5PHIA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D5PHIA_wea,
        addra     => FM_BBBB_D5PHIA_writeaddr,
        dina      => FM_BBBB_D5PHIA_din,
        wea_out       => FM_BBBB_D5PHIA_wea_delay,
        addra_out     => FM_BBBB_D5PHIA_writeaddr_delay,
        dina_out      => FM_BBBB_D5PHIA_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D5PHIA_start
      );

    FM_AAAA_D5PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D5PHIB_wea_delay,
        addra     => FM_AAAA_D5PHIB_writeaddr_delay,
        dina      => FM_AAAA_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D5PHIB_V_readaddr,
        doutb     => FM_AAAA_D5PHIB_V_dout,
        sync_nent => FM_AAAA_D5PHIB_start,
        nent_o    => FM_AAAA_D5PHIB_AV_dout_nent
      );

    FM_AAAA_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D5PHIB_wea,
        addra     => FM_AAAA_D5PHIB_writeaddr,
        dina      => FM_AAAA_D5PHIB_din,
        wea_out       => FM_AAAA_D5PHIB_wea_delay,
        addra_out     => FM_AAAA_D5PHIB_writeaddr_delay,
        dina_out      => FM_AAAA_D5PHIB_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D5PHIB_start
      );

    FM_BBBB_D5PHIB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D5PHIB"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D5PHIB_wea_delay,
        addra     => FM_BBBB_D5PHIB_writeaddr_delay,
        dina      => FM_BBBB_D5PHIB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D5PHIB_V_readaddr,
        doutb     => FM_BBBB_D5PHIB_V_dout,
        sync_nent => FM_BBBB_D5PHIB_start,
        nent_o    => FM_BBBB_D5PHIB_AV_dout_nent
      );

    FM_BBBB_D5PHIB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D5PHIB_wea,
        addra     => FM_BBBB_D5PHIB_writeaddr,
        dina      => FM_BBBB_D5PHIB_din,
        wea_out       => FM_BBBB_D5PHIB_wea_delay,
        addra_out     => FM_BBBB_D5PHIB_writeaddr_delay,
        dina_out      => FM_BBBB_D5PHIB_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D5PHIB_start
      );

    FM_AAAA_D5PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D5PHIC_wea_delay,
        addra     => FM_AAAA_D5PHIC_writeaddr_delay,
        dina      => FM_AAAA_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D5PHIC_V_readaddr,
        doutb     => FM_AAAA_D5PHIC_V_dout,
        sync_nent => FM_AAAA_D5PHIC_start,
        nent_o    => FM_AAAA_D5PHIC_AV_dout_nent
      );

    FM_AAAA_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D5PHIC_wea,
        addra     => FM_AAAA_D5PHIC_writeaddr,
        dina      => FM_AAAA_D5PHIC_din,
        wea_out       => FM_AAAA_D5PHIC_wea_delay,
        addra_out     => FM_AAAA_D5PHIC_writeaddr_delay,
        dina_out      => FM_AAAA_D5PHIC_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D5PHIC_start
      );

    FM_BBBB_D5PHIC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D5PHIC"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D5PHIC_wea_delay,
        addra     => FM_BBBB_D5PHIC_writeaddr_delay,
        dina      => FM_BBBB_D5PHIC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D5PHIC_V_readaddr,
        doutb     => FM_BBBB_D5PHIC_V_dout,
        sync_nent => FM_BBBB_D5PHIC_start,
        nent_o    => FM_BBBB_D5PHIC_AV_dout_nent
      );

    FM_BBBB_D5PHIC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D5PHIC_wea,
        addra     => FM_BBBB_D5PHIC_writeaddr,
        dina      => FM_BBBB_D5PHIC_din,
        wea_out       => FM_BBBB_D5PHIC_wea_delay,
        addra_out     => FM_BBBB_D5PHIC_writeaddr_delay,
        dina_out      => FM_BBBB_D5PHIC_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D5PHIC_start
      );

    FM_AAAA_D5PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_AAAA_D5PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_AAAA_D5PHID_wea_delay,
        addra     => FM_AAAA_D5PHID_writeaddr_delay,
        dina      => FM_AAAA_D5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_AAAA_D5PHID_V_readaddr,
        doutb     => FM_AAAA_D5PHID_V_dout,
        sync_nent => FM_AAAA_D5PHID_start,
        nent_o    => FM_AAAA_D5PHID_AV_dout_nent
      );

    FM_AAAA_D5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_AAAA_D5PHID_wea,
        addra     => FM_AAAA_D5PHID_writeaddr,
        dina      => FM_AAAA_D5PHID_din,
        wea_out       => FM_AAAA_D5PHID_wea_delay,
        addra_out     => FM_AAAA_D5PHID_writeaddr_delay,
        dina_out      => FM_AAAA_D5PHID_din_delay,
        done       => MP_done,
        start      => FM_AAAA_D5PHID_start
      );

    FM_BBBB_D5PHID : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 55,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "FM_BBBB_D5PHID"
      )
      port map (
        clka      => clk,
        wea       => FM_BBBB_D5PHID_wea_delay,
        addra     => FM_BBBB_D5PHID_writeaddr_delay,
        dina      => FM_BBBB_D5PHID_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => FM_BBBB_D5PHID_V_readaddr,
        doutb     => FM_BBBB_D5PHID_V_dout,
        sync_nent => FM_BBBB_D5PHID_start,
        nent_o    => FM_BBBB_D5PHID_AV_dout_nent
      );

    FM_BBBB_D5PHID_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 55
      )
      port map (
        clk      => clk,
        wea       => FM_BBBB_D5PHID_wea,
        addra     => FM_BBBB_D5PHID_writeaddr,
        dina      => FM_BBBB_D5PHID_din,
        wea_out       => FM_BBBB_D5PHID_wea_delay,
        addra_out     => FM_BBBB_D5PHID_writeaddr_delay,
        dina_out      => FM_BBBB_D5PHID_din_delay,
        done       => MP_done,
        start      => FM_BBBB_D5PHID_start
      );

  VMSMER_L1PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIA_bx_in,
      start => VMSMER_L1PHIA_start,
      enb   => AS_L1PHIAin_enb,
      addra => AS_L1PHIAin_V_readaddr,
      din   => AS_L1PHIAin_V_dout,
      dout  => AS_L1PHIAin_V_as,
      valid  => AS_L1PHIAin_valid,
      index  => AS_L1PHIAin_index(6 downto 0),
      nent  => AS_L1PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIA_bx_in,
      start => VMSMER_L1PHIA_start
  );

  LATCH_VMSMER_L1PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIA_bx
  );

  VMSMER_L1PHIA : entity work.VMSMER_L1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIA_bx,
      valid        => AS_L1PHIAin_valid,
      index        => AS_L1PHIAin_index,
      allStub_data_V        => AS_L1PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIAn2_din
  );

  VMSMER_L1PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIB_bx_in,
      start => VMSMER_L1PHIB_start,
      enb   => AS_L1PHIBin_enb,
      addra => AS_L1PHIBin_V_readaddr,
      din   => AS_L1PHIBin_V_dout,
      dout  => AS_L1PHIBin_V_as,
      valid  => AS_L1PHIBin_valid,
      index  => AS_L1PHIBin_index(6 downto 0),
      nent  => AS_L1PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIB_bx_in,
      start => VMSMER_L1PHIB_start
  );

  LATCH_VMSMER_L1PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIB_bx
  );

  VMSMER_L1PHIB : entity work.VMSMER_L1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIB_bx,
      valid        => AS_L1PHIBin_valid,
      index        => AS_L1PHIBin_index,
      allStub_data_V        => AS_L1PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIBn2_din
  );

  VMSMER_L1PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIC_bx_in,
      start => VMSMER_L1PHIC_start,
      enb   => AS_L1PHICin_enb,
      addra => AS_L1PHICin_V_readaddr,
      din   => AS_L1PHICin_V_dout,
      dout  => AS_L1PHICin_V_as,
      valid  => AS_L1PHICin_valid,
      index  => AS_L1PHICin_index(6 downto 0),
      nent  => AS_L1PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIC_bx_in,
      start => VMSMER_L1PHIC_start
  );

  LATCH_VMSMER_L1PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIC_bx
  );

  VMSMER_L1PHIC : entity work.VMSMER_L1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIC_bx,
      valid        => AS_L1PHICin_valid,
      index        => AS_L1PHICin_index,
      allStub_data_V        => AS_L1PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHICn2_din
  );

  VMSMER_L1PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHID_bx_in,
      start => VMSMER_L1PHID_start,
      enb   => AS_L1PHIDin_enb,
      addra => AS_L1PHIDin_V_readaddr,
      din   => AS_L1PHIDin_V_dout,
      dout  => AS_L1PHIDin_V_as,
      valid  => AS_L1PHIDin_valid,
      index  => AS_L1PHIDin_index(6 downto 0),
      nent  => AS_L1PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHID_bx_in,
      start => VMSMER_L1PHID_start
  );

  LATCH_VMSMER_L1PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHID_bx
  );

  VMSMER_L1PHID : entity work.VMSMER_L1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHID_bx,
      valid        => AS_L1PHIDin_valid,
      index        => AS_L1PHIDin_index,
      allStub_data_V        => AS_L1PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIDn2_din
  );

  VMSMER_L1PHIE_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIE_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIE_bx_in,
      start => VMSMER_L1PHIE_start,
      enb   => AS_L1PHIEin_enb,
      addra => AS_L1PHIEin_V_readaddr,
      din   => AS_L1PHIEin_V_dout,
      dout  => AS_L1PHIEin_V_as,
      valid  => AS_L1PHIEin_valid,
      index  => AS_L1PHIEin_index(6 downto 0),
      nent  => AS_L1PHIEin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIE: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIE_bx_in,
      start => VMSMER_L1PHIE_start
  );

  LATCH_VMSMER_L1PHIE_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIE_bx
  );

  VMSMER_L1PHIE : entity work.VMSMER_L1PHIE
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIE_bx,
      valid        => AS_L1PHIEin_valid,
      index        => AS_L1PHIEin_index,
      allStub_data_V        => AS_L1PHIEin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIEn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIEn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIEn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIEn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIEn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIEn2_din
  );

  VMSMER_L1PHIF_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIF_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIF_bx_in,
      start => VMSMER_L1PHIF_start,
      enb   => AS_L1PHIFin_enb,
      addra => AS_L1PHIFin_V_readaddr,
      din   => AS_L1PHIFin_V_dout,
      dout  => AS_L1PHIFin_V_as,
      valid  => AS_L1PHIFin_valid,
      index  => AS_L1PHIFin_index(6 downto 0),
      nent  => AS_L1PHIFin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIF: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIF_bx_in,
      start => VMSMER_L1PHIF_start
  );

  LATCH_VMSMER_L1PHIF_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIF_bx
  );

  VMSMER_L1PHIF : entity work.VMSMER_L1PHIF
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIF_bx,
      valid        => AS_L1PHIFin_valid,
      index        => AS_L1PHIFin_index,
      allStub_data_V        => AS_L1PHIFin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIFn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIFn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIFn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIFn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIFn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIFn2_din
  );

  VMSMER_L1PHIG_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIG_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIG_bx_in,
      start => VMSMER_L1PHIG_start,
      enb   => AS_L1PHIGin_enb,
      addra => AS_L1PHIGin_V_readaddr,
      din   => AS_L1PHIGin_V_dout,
      dout  => AS_L1PHIGin_V_as,
      valid  => AS_L1PHIGin_valid,
      index  => AS_L1PHIGin_index(6 downto 0),
      nent  => AS_L1PHIGin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIG: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIG_bx_in,
      start => VMSMER_L1PHIG_start
  );

  LATCH_VMSMER_L1PHIG_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIG_bx
  );

  VMSMER_L1PHIG : entity work.VMSMER_L1PHIG
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIG_bx,
      valid        => AS_L1PHIGin_valid,
      index        => AS_L1PHIGin_index,
      allStub_data_V        => AS_L1PHIGin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIGn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIGn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIGn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIGn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIGn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIGn2_din
  );

  VMSMER_L1PHIH_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L1PHIH_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L1PHIH_bx_in,
      start => VMSMER_L1PHIH_start,
      enb   => AS_L1PHIHin_enb,
      addra => AS_L1PHIHin_V_readaddr,
      din   => AS_L1PHIHin_V_dout,
      dout  => AS_L1PHIHin_V_as,
      valid  => AS_L1PHIHin_valid,
      index  => AS_L1PHIHin_index(6 downto 0),
      nent  => AS_L1PHIHin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L1PHIH: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIH_bx_in,
      start => VMSMER_L1PHIH_start
  );

  LATCH_VMSMER_L1PHIH_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L1PHIH_bx
  );

  VMSMER_L1PHIH : entity work.VMSMER_L1PHIH
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L1PHIH_bx,
      valid        => AS_L1PHIHin_valid,
      index        => AS_L1PHIHin_index,
      allStub_data_V        => AS_L1PHIHin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L1PHIHn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L1PHIHn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L1PHIHn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIHn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIHn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIHn2_din
  );

  VMSMER_L2PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L2PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L2PHIA_bx_in,
      start => VMSMER_L2PHIA_start,
      enb   => AS_L2PHIAin_enb,
      addra => AS_L2PHIAin_V_readaddr,
      din   => AS_L2PHIAin_V_dout,
      dout  => AS_L2PHIAin_V_as,
      valid  => AS_L2PHIAin_valid,
      index  => AS_L2PHIAin_index(6 downto 0),
      nent  => AS_L2PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIA_bx_in,
      start => VMSMER_L2PHIA_start
  );

  LATCH_VMSMER_L2PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIA_bx
  );

  VMSMER_L2PHIA : entity work.VMSMER_L2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L2PHIA_bx,
      valid        => AS_L2PHIAin_valid,
      index        => AS_L2PHIAin_index,
      allStub_data_V        => AS_L2PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L2PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L2PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L2PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIAn2_din
  );

  VMSMER_L2PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L2PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L2PHIB_bx_in,
      start => VMSMER_L2PHIB_start,
      enb   => AS_L2PHIBin_enb,
      addra => AS_L2PHIBin_V_readaddr,
      din   => AS_L2PHIBin_V_dout,
      dout  => AS_L2PHIBin_V_as,
      valid  => AS_L2PHIBin_valid,
      index  => AS_L2PHIBin_index(6 downto 0),
      nent  => AS_L2PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIB_bx_in,
      start => VMSMER_L2PHIB_start
  );

  LATCH_VMSMER_L2PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIB_bx
  );

  VMSMER_L2PHIB : entity work.VMSMER_L2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L2PHIB_bx,
      valid        => AS_L2PHIBin_valid,
      index        => AS_L2PHIBin_index,
      allStub_data_V        => AS_L2PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L2PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L2PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L2PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIBn2_din
  );

  VMSMER_L2PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L2PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L2PHIC_bx_in,
      start => VMSMER_L2PHIC_start,
      enb   => AS_L2PHICin_enb,
      addra => AS_L2PHICin_V_readaddr,
      din   => AS_L2PHICin_V_dout,
      dout  => AS_L2PHICin_V_as,
      valid  => AS_L2PHICin_valid,
      index  => AS_L2PHICin_index(6 downto 0),
      nent  => AS_L2PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIC_bx_in,
      start => VMSMER_L2PHIC_start
  );

  LATCH_VMSMER_L2PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHIC_bx
  );

  VMSMER_L2PHIC : entity work.VMSMER_L2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L2PHIC_bx,
      valid        => AS_L2PHICin_valid,
      index        => AS_L2PHICin_index,
      allStub_data_V        => AS_L2PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L2PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L2PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L2PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHICn2_din
  );

  VMSMER_L2PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L2PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L2PHID_bx_in,
      start => VMSMER_L2PHID_start,
      enb   => AS_L2PHIDin_enb,
      addra => AS_L2PHIDin_V_readaddr,
      din   => AS_L2PHIDin_V_dout,
      dout  => AS_L2PHIDin_V_as,
      valid  => AS_L2PHIDin_valid,
      index  => AS_L2PHIDin_index(6 downto 0),
      nent  => AS_L2PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHID_bx_in,
      start => VMSMER_L2PHID_start
  );

  LATCH_VMSMER_L2PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L2PHID_bx
  );

  VMSMER_L2PHID : entity work.VMSMER_L2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L2PHID_bx,
      valid        => AS_L2PHIDin_valid,
      index        => AS_L2PHIDin_index,
      allStub_data_V        => AS_L2PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L2PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L2PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L2PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIDn2_din
  );

  VMSMER_L3PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L3PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L3PHIA_bx_in,
      start => VMSMER_L3PHIA_start,
      enb   => AS_L3PHIAin_enb,
      addra => AS_L3PHIAin_V_readaddr,
      din   => AS_L3PHIAin_V_dout,
      dout  => AS_L3PHIAin_V_as,
      valid  => AS_L3PHIAin_valid,
      index  => AS_L3PHIAin_index(6 downto 0),
      nent  => AS_L3PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIA_bx_in,
      start => VMSMER_L3PHIA_start
  );

  LATCH_VMSMER_L3PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIA_bx
  );

  VMSMER_L3PHIA : entity work.VMSMER_L3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L3PHIA_bx,
      valid        => AS_L3PHIAin_valid,
      index        => AS_L3PHIAin_index,
      allStub_data_V        => AS_L3PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L3PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L3PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L3PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIAn2_din
  );

  VMSMER_L3PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L3PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L3PHIB_bx_in,
      start => VMSMER_L3PHIB_start,
      enb   => AS_L3PHIBin_enb,
      addra => AS_L3PHIBin_V_readaddr,
      din   => AS_L3PHIBin_V_dout,
      dout  => AS_L3PHIBin_V_as,
      valid  => AS_L3PHIBin_valid,
      index  => AS_L3PHIBin_index(6 downto 0),
      nent  => AS_L3PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIB_bx_in,
      start => VMSMER_L3PHIB_start
  );

  LATCH_VMSMER_L3PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIB_bx
  );

  VMSMER_L3PHIB : entity work.VMSMER_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L3PHIB_bx,
      valid        => AS_L3PHIBin_valid,
      index        => AS_L3PHIBin_index,
      allStub_data_V        => AS_L3PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L3PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L3PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L3PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIBn2_din
  );

  VMSMER_L3PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L3PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L3PHIC_bx_in,
      start => VMSMER_L3PHIC_start,
      enb   => AS_L3PHICin_enb,
      addra => AS_L3PHICin_V_readaddr,
      din   => AS_L3PHICin_V_dout,
      dout  => AS_L3PHICin_V_as,
      valid  => AS_L3PHICin_valid,
      index  => AS_L3PHICin_index(6 downto 0),
      nent  => AS_L3PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIC_bx_in,
      start => VMSMER_L3PHIC_start
  );

  LATCH_VMSMER_L3PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHIC_bx
  );

  VMSMER_L3PHIC : entity work.VMSMER_L3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L3PHIC_bx,
      valid        => AS_L3PHICin_valid,
      index        => AS_L3PHICin_index,
      allStub_data_V        => AS_L3PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L3PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L3PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L3PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHICn2_din
  );

  VMSMER_L3PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L3PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L3PHID_bx_in,
      start => VMSMER_L3PHID_start,
      enb   => AS_L3PHIDin_enb,
      addra => AS_L3PHIDin_V_readaddr,
      din   => AS_L3PHIDin_V_dout,
      dout  => AS_L3PHIDin_V_as,
      valid  => AS_L3PHIDin_valid,
      index  => AS_L3PHIDin_index(6 downto 0),
      nent  => AS_L3PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHID_bx_in,
      start => VMSMER_L3PHID_start
  );

  LATCH_VMSMER_L3PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L3PHID_bx
  );

  VMSMER_L3PHID : entity work.VMSMER_L3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L3PHID_bx,
      valid        => AS_L3PHIDin_valid,
      index        => AS_L3PHIDin_index,
      allStub_data_V        => AS_L3PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L3PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L3PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L3PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIDn2_din
  );

  VMSMER_L4PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L4PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L4PHIA_bx_in,
      start => VMSMER_L4PHIA_start,
      enb   => AS_L4PHIAin_enb,
      addra => AS_L4PHIAin_V_readaddr,
      din   => AS_L4PHIAin_V_dout,
      dout  => AS_L4PHIAin_V_as,
      valid  => AS_L4PHIAin_valid,
      index  => AS_L4PHIAin_index(6 downto 0),
      nent  => AS_L4PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIA_bx_in,
      start => VMSMER_L4PHIA_start
  );

  LATCH_VMSMER_L4PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIA_bx
  );

  VMSMER_L4PHIA : entity work.VMSMER_L4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L4PHIA_bx,
      valid        => AS_L4PHIAin_valid,
      index        => AS_L4PHIAin_index,
      allStub_data_V        => AS_L4PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L4PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L4PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L4PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIAn2_din
  );

  VMSMER_L4PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L4PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L4PHIB_bx_in,
      start => VMSMER_L4PHIB_start,
      enb   => AS_L4PHIBin_enb,
      addra => AS_L4PHIBin_V_readaddr,
      din   => AS_L4PHIBin_V_dout,
      dout  => AS_L4PHIBin_V_as,
      valid  => AS_L4PHIBin_valid,
      index  => AS_L4PHIBin_index(6 downto 0),
      nent  => AS_L4PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIB_bx_in,
      start => VMSMER_L4PHIB_start
  );

  LATCH_VMSMER_L4PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIB_bx
  );

  VMSMER_L4PHIB : entity work.VMSMER_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L4PHIB_bx,
      valid        => AS_L4PHIBin_valid,
      index        => AS_L4PHIBin_index,
      allStub_data_V        => AS_L4PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L4PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L4PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L4PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIBn2_din
  );

  VMSMER_L4PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L4PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L4PHIC_bx_in,
      start => VMSMER_L4PHIC_start,
      enb   => AS_L4PHICin_enb,
      addra => AS_L4PHICin_V_readaddr,
      din   => AS_L4PHICin_V_dout,
      dout  => AS_L4PHICin_V_as,
      valid  => AS_L4PHICin_valid,
      index  => AS_L4PHICin_index(6 downto 0),
      nent  => AS_L4PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIC_bx_in,
      start => VMSMER_L4PHIC_start
  );

  LATCH_VMSMER_L4PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHIC_bx
  );

  VMSMER_L4PHIC : entity work.VMSMER_L4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L4PHIC_bx,
      valid        => AS_L4PHICin_valid,
      index        => AS_L4PHICin_index,
      allStub_data_V        => AS_L4PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L4PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L4PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L4PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHICn2_din
  );

  VMSMER_L4PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L4PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L4PHID_bx_in,
      start => VMSMER_L4PHID_start,
      enb   => AS_L4PHIDin_enb,
      addra => AS_L4PHIDin_V_readaddr,
      din   => AS_L4PHIDin_V_dout,
      dout  => AS_L4PHIDin_V_as,
      valid  => AS_L4PHIDin_valid,
      index  => AS_L4PHIDin_index(6 downto 0),
      nent  => AS_L4PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHID_bx_in,
      start => VMSMER_L4PHID_start
  );

  LATCH_VMSMER_L4PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L4PHID_bx
  );

  VMSMER_L4PHID : entity work.VMSMER_L4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L4PHID_bx,
      valid        => AS_L4PHIDin_valid,
      index        => AS_L4PHIDin_index,
      allStub_data_V        => AS_L4PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L4PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L4PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L4PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIDn2_din
  );

  VMSMER_L5PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L5PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L5PHIA_bx_in,
      start => VMSMER_L5PHIA_start,
      enb   => AS_L5PHIAin_enb,
      addra => AS_L5PHIAin_V_readaddr,
      din   => AS_L5PHIAin_V_dout,
      dout  => AS_L5PHIAin_V_as,
      valid  => AS_L5PHIAin_valid,
      index  => AS_L5PHIAin_index(6 downto 0),
      nent  => AS_L5PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIA_bx_in,
      start => VMSMER_L5PHIA_start
  );

  LATCH_VMSMER_L5PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIA_bx
  );

  VMSMER_L5PHIA : entity work.VMSMER_L5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L5PHIA_bx,
      valid        => AS_L5PHIAin_valid,
      index        => AS_L5PHIAin_index,
      allStub_data_V        => AS_L5PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L5PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L5PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L5PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIAn2_din
  );

  VMSMER_L5PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L5PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L5PHIB_bx_in,
      start => VMSMER_L5PHIB_start,
      enb   => AS_L5PHIBin_enb,
      addra => AS_L5PHIBin_V_readaddr,
      din   => AS_L5PHIBin_V_dout,
      dout  => AS_L5PHIBin_V_as,
      valid  => AS_L5PHIBin_valid,
      index  => AS_L5PHIBin_index(6 downto 0),
      nent  => AS_L5PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIB_bx_in,
      start => VMSMER_L5PHIB_start
  );

  LATCH_VMSMER_L5PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIB_bx
  );

  VMSMER_L5PHIB : entity work.VMSMER_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L5PHIB_bx,
      valid        => AS_L5PHIBin_valid,
      index        => AS_L5PHIBin_index,
      allStub_data_V        => AS_L5PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L5PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L5PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L5PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIBn2_din
  );

  VMSMER_L5PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L5PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L5PHIC_bx_in,
      start => VMSMER_L5PHIC_start,
      enb   => AS_L5PHICin_enb,
      addra => AS_L5PHICin_V_readaddr,
      din   => AS_L5PHICin_V_dout,
      dout  => AS_L5PHICin_V_as,
      valid  => AS_L5PHICin_valid,
      index  => AS_L5PHICin_index(6 downto 0),
      nent  => AS_L5PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIC_bx_in,
      start => VMSMER_L5PHIC_start
  );

  LATCH_VMSMER_L5PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHIC_bx
  );

  VMSMER_L5PHIC : entity work.VMSMER_L5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L5PHIC_bx,
      valid        => AS_L5PHICin_valid,
      index        => AS_L5PHICin_index,
      allStub_data_V        => AS_L5PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L5PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L5PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L5PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHICn2_din
  );

  VMSMER_L5PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L5PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L5PHID_bx_in,
      start => VMSMER_L5PHID_start,
      enb   => AS_L5PHIDin_enb,
      addra => AS_L5PHIDin_V_readaddr,
      din   => AS_L5PHIDin_V_dout,
      dout  => AS_L5PHIDin_V_as,
      valid  => AS_L5PHIDin_valid,
      index  => AS_L5PHIDin_index(6 downto 0),
      nent  => AS_L5PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHID_bx_in,
      start => VMSMER_L5PHID_start
  );

  LATCH_VMSMER_L5PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L5PHID_bx
  );

  VMSMER_L5PHID : entity work.VMSMER_L5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L5PHID_bx,
      valid        => AS_L5PHIDin_valid,
      index        => AS_L5PHIDin_index,
      allStub_data_V        => AS_L5PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L5PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L5PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L5PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIDn2_din
  );

  VMSMER_L6PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L6PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L6PHIA_bx_in,
      start => VMSMER_L6PHIA_start,
      enb   => AS_L6PHIAin_enb,
      addra => AS_L6PHIAin_V_readaddr,
      din   => AS_L6PHIAin_V_dout,
      dout  => AS_L6PHIAin_V_as,
      valid  => AS_L6PHIAin_valid,
      index  => AS_L6PHIAin_index(6 downto 0),
      nent  => AS_L6PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L6PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIA_bx_in,
      start => VMSMER_L6PHIA_start
  );

  LATCH_VMSMER_L6PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIA_bx
  );

  VMSMER_L6PHIA : entity work.VMSMER_L6PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L6PHIA_bx,
      valid        => AS_L6PHIAin_valid,
      index        => AS_L6PHIAin_index,
      allStub_data_V        => AS_L6PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L6PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L6PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L6PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIAn2_din
  );

  VMSMER_L6PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L6PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L6PHIB_bx_in,
      start => VMSMER_L6PHIB_start,
      enb   => AS_L6PHIBin_enb,
      addra => AS_L6PHIBin_V_readaddr,
      din   => AS_L6PHIBin_V_dout,
      dout  => AS_L6PHIBin_V_as,
      valid  => AS_L6PHIBin_valid,
      index  => AS_L6PHIBin_index(6 downto 0),
      nent  => AS_L6PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L6PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIB_bx_in,
      start => VMSMER_L6PHIB_start
  );

  LATCH_VMSMER_L6PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIB_bx
  );

  VMSMER_L6PHIB : entity work.VMSMER_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L6PHIB_bx,
      valid        => AS_L6PHIBin_valid,
      index        => AS_L6PHIBin_index,
      allStub_data_V        => AS_L6PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L6PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L6PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L6PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIBn2_din
  );

  VMSMER_L6PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L6PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L6PHIC_bx_in,
      start => VMSMER_L6PHIC_start,
      enb   => AS_L6PHICin_enb,
      addra => AS_L6PHICin_V_readaddr,
      din   => AS_L6PHICin_V_dout,
      dout  => AS_L6PHICin_V_as,
      valid  => AS_L6PHICin_valid,
      index  => AS_L6PHICin_index(6 downto 0),
      nent  => AS_L6PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L6PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIC_bx_in,
      start => VMSMER_L6PHIC_start
  );

  LATCH_VMSMER_L6PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHIC_bx
  );

  VMSMER_L6PHIC : entity work.VMSMER_L6PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L6PHIC_bx,
      valid        => AS_L6PHICin_valid,
      index        => AS_L6PHICin_index,
      allStub_data_V        => AS_L6PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L6PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L6PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L6PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHICn2_din
  );

  VMSMER_L6PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_L6PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_L6PHID_bx_in,
      start => VMSMER_L6PHID_start,
      enb   => AS_L6PHIDin_enb,
      addra => AS_L6PHIDin_V_readaddr,
      din   => AS_L6PHIDin_V_dout,
      dout  => AS_L6PHIDin_V_as,
      valid  => AS_L6PHIDin_valid,
      index  => AS_L6PHIDin_index(6 downto 0),
      nent  => AS_L6PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_L6PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHID_bx_in,
      start => VMSMER_L6PHID_start
  );

  LATCH_VMSMER_L6PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_L6PHID_bx
  );

  VMSMER_L6PHID : entity work.VMSMER_L6PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_L6PHID_bx,
      valid        => AS_L6PHIDin_valid,
      index        => AS_L6PHIDin_index,
      allStub_data_V        => AS_L6PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_L6PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_L6PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_L6PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIDn2_din
  );

  VMSMER_D1PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D1PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D1PHIA_bx_in,
      start => VMSMER_D1PHIA_start,
      enb   => AS_D1PHIAin_enb,
      addra => AS_D1PHIAin_V_readaddr,
      din   => AS_D1PHIAin_V_dout,
      dout  => AS_D1PHIAin_V_as,
      valid  => AS_D1PHIAin_valid,
      index  => AS_D1PHIAin_index(6 downto 0),
      nent  => AS_D1PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIA_bx_in,
      start => VMSMER_D1PHIA_start
  );

  LATCH_VMSMER_D1PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIA_bx
  );

  VMSMER_D1PHIA : entity work.VMSMER_D1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D1PHIA_bx,
      valid        => AS_D1PHIAin_valid,
      index        => AS_D1PHIAin_index,
      allStub_data_V        => AS_D1PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D1PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D1PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D1PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIAn2_din
  );

  VMSMER_D1PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D1PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D1PHIB_bx_in,
      start => VMSMER_D1PHIB_start,
      enb   => AS_D1PHIBin_enb,
      addra => AS_D1PHIBin_V_readaddr,
      din   => AS_D1PHIBin_V_dout,
      dout  => AS_D1PHIBin_V_as,
      valid  => AS_D1PHIBin_valid,
      index  => AS_D1PHIBin_index(6 downto 0),
      nent  => AS_D1PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIB_bx_in,
      start => VMSMER_D1PHIB_start
  );

  LATCH_VMSMER_D1PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIB_bx
  );

  VMSMER_D1PHIB : entity work.VMSMER_D1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D1PHIB_bx,
      valid        => AS_D1PHIBin_valid,
      index        => AS_D1PHIBin_index,
      allStub_data_V        => AS_D1PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D1PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D1PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D1PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIBn2_din
  );

  VMSMER_D1PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D1PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D1PHIC_bx_in,
      start => VMSMER_D1PHIC_start,
      enb   => AS_D1PHICin_enb,
      addra => AS_D1PHICin_V_readaddr,
      din   => AS_D1PHICin_V_dout,
      dout  => AS_D1PHICin_V_as,
      valid  => AS_D1PHICin_valid,
      index  => AS_D1PHICin_index(6 downto 0),
      nent  => AS_D1PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIC_bx_in,
      start => VMSMER_D1PHIC_start
  );

  LATCH_VMSMER_D1PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHIC_bx
  );

  VMSMER_D1PHIC : entity work.VMSMER_D1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D1PHIC_bx,
      valid        => AS_D1PHICin_valid,
      index        => AS_D1PHICin_index,
      allStub_data_V        => AS_D1PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D1PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D1PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D1PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHICn2_din
  );

  VMSMER_D1PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D1PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D1PHID_bx_in,
      start => VMSMER_D1PHID_start,
      enb   => AS_D1PHIDin_enb,
      addra => AS_D1PHIDin_V_readaddr,
      din   => AS_D1PHIDin_V_dout,
      dout  => AS_D1PHIDin_V_as,
      valid  => AS_D1PHIDin_valid,
      index  => AS_D1PHIDin_index(6 downto 0),
      nent  => AS_D1PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHID_bx_in,
      start => VMSMER_D1PHID_start
  );

  LATCH_VMSMER_D1PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D1PHID_bx
  );

  VMSMER_D1PHID : entity work.VMSMER_D1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D1PHID_bx,
      valid        => AS_D1PHIDin_valid,
      index        => AS_D1PHIDin_index,
      allStub_data_V        => AS_D1PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D1PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D1PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D1PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIDn2_din
  );

  VMSMER_D2PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D2PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D2PHIA_bx_in,
      start => VMSMER_D2PHIA_start,
      enb   => AS_D2PHIAin_enb,
      addra => AS_D2PHIAin_V_readaddr,
      din   => AS_D2PHIAin_V_dout,
      dout  => AS_D2PHIAin_V_as,
      valid  => AS_D2PHIAin_valid,
      index  => AS_D2PHIAin_index(6 downto 0),
      nent  => AS_D2PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIA_bx_in,
      start => VMSMER_D2PHIA_start
  );

  LATCH_VMSMER_D2PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIA_bx
  );

  VMSMER_D2PHIA : entity work.VMSMER_D2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D2PHIA_bx,
      valid        => AS_D2PHIAin_valid,
      index        => AS_D2PHIAin_index,
      allStub_data_V        => AS_D2PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D2PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D2PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D2PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIAn2_din
  );

  VMSMER_D2PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D2PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D2PHIB_bx_in,
      start => VMSMER_D2PHIB_start,
      enb   => AS_D2PHIBin_enb,
      addra => AS_D2PHIBin_V_readaddr,
      din   => AS_D2PHIBin_V_dout,
      dout  => AS_D2PHIBin_V_as,
      valid  => AS_D2PHIBin_valid,
      index  => AS_D2PHIBin_index(6 downto 0),
      nent  => AS_D2PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIB_bx_in,
      start => VMSMER_D2PHIB_start
  );

  LATCH_VMSMER_D2PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIB_bx
  );

  VMSMER_D2PHIB : entity work.VMSMER_D2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D2PHIB_bx,
      valid        => AS_D2PHIBin_valid,
      index        => AS_D2PHIBin_index,
      allStub_data_V        => AS_D2PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D2PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D2PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D2PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIBn2_din
  );

  VMSMER_D2PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D2PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D2PHIC_bx_in,
      start => VMSMER_D2PHIC_start,
      enb   => AS_D2PHICin_enb,
      addra => AS_D2PHICin_V_readaddr,
      din   => AS_D2PHICin_V_dout,
      dout  => AS_D2PHICin_V_as,
      valid  => AS_D2PHICin_valid,
      index  => AS_D2PHICin_index(6 downto 0),
      nent  => AS_D2PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIC_bx_in,
      start => VMSMER_D2PHIC_start
  );

  LATCH_VMSMER_D2PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHIC_bx
  );

  VMSMER_D2PHIC : entity work.VMSMER_D2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D2PHIC_bx,
      valid        => AS_D2PHICin_valid,
      index        => AS_D2PHICin_index,
      allStub_data_V        => AS_D2PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D2PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D2PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D2PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHICn2_din
  );

  VMSMER_D2PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D2PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D2PHID_bx_in,
      start => VMSMER_D2PHID_start,
      enb   => AS_D2PHIDin_enb,
      addra => AS_D2PHIDin_V_readaddr,
      din   => AS_D2PHIDin_V_dout,
      dout  => AS_D2PHIDin_V_as,
      valid  => AS_D2PHIDin_valid,
      index  => AS_D2PHIDin_index(6 downto 0),
      nent  => AS_D2PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHID_bx_in,
      start => VMSMER_D2PHID_start
  );

  LATCH_VMSMER_D2PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D2PHID_bx
  );

  VMSMER_D2PHID : entity work.VMSMER_D2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D2PHID_bx,
      valid        => AS_D2PHIDin_valid,
      index        => AS_D2PHIDin_index,
      allStub_data_V        => AS_D2PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D2PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D2PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D2PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIDn2_din
  );

  VMSMER_D3PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D3PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D3PHIA_bx_in,
      start => VMSMER_D3PHIA_start,
      enb   => AS_D3PHIAin_enb,
      addra => AS_D3PHIAin_V_readaddr,
      din   => AS_D3PHIAin_V_dout,
      dout  => AS_D3PHIAin_V_as,
      valid  => AS_D3PHIAin_valid,
      index  => AS_D3PHIAin_index(6 downto 0),
      nent  => AS_D3PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIA_bx_in,
      start => VMSMER_D3PHIA_start
  );

  LATCH_VMSMER_D3PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIA_bx
  );

  VMSMER_D3PHIA : entity work.VMSMER_D3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D3PHIA_bx,
      valid        => AS_D3PHIAin_valid,
      index        => AS_D3PHIAin_index,
      allStub_data_V        => AS_D3PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D3PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D3PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D3PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIAn2_din
  );

  VMSMER_D3PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D3PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D3PHIB_bx_in,
      start => VMSMER_D3PHIB_start,
      enb   => AS_D3PHIBin_enb,
      addra => AS_D3PHIBin_V_readaddr,
      din   => AS_D3PHIBin_V_dout,
      dout  => AS_D3PHIBin_V_as,
      valid  => AS_D3PHIBin_valid,
      index  => AS_D3PHIBin_index(6 downto 0),
      nent  => AS_D3PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIB_bx_in,
      start => VMSMER_D3PHIB_start
  );

  LATCH_VMSMER_D3PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIB_bx
  );

  VMSMER_D3PHIB : entity work.VMSMER_D3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D3PHIB_bx,
      valid        => AS_D3PHIBin_valid,
      index        => AS_D3PHIBin_index,
      allStub_data_V        => AS_D3PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D3PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D3PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D3PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIBn2_din
  );

  VMSMER_D3PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D3PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D3PHIC_bx_in,
      start => VMSMER_D3PHIC_start,
      enb   => AS_D3PHICin_enb,
      addra => AS_D3PHICin_V_readaddr,
      din   => AS_D3PHICin_V_dout,
      dout  => AS_D3PHICin_V_as,
      valid  => AS_D3PHICin_valid,
      index  => AS_D3PHICin_index(6 downto 0),
      nent  => AS_D3PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIC_bx_in,
      start => VMSMER_D3PHIC_start
  );

  LATCH_VMSMER_D3PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHIC_bx
  );

  VMSMER_D3PHIC : entity work.VMSMER_D3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D3PHIC_bx,
      valid        => AS_D3PHICin_valid,
      index        => AS_D3PHICin_index,
      allStub_data_V        => AS_D3PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D3PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D3PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D3PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHICn2_din
  );

  VMSMER_D3PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D3PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D3PHID_bx_in,
      start => VMSMER_D3PHID_start,
      enb   => AS_D3PHIDin_enb,
      addra => AS_D3PHIDin_V_readaddr,
      din   => AS_D3PHIDin_V_dout,
      dout  => AS_D3PHIDin_V_as,
      valid  => AS_D3PHIDin_valid,
      index  => AS_D3PHIDin_index(6 downto 0),
      nent  => AS_D3PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHID_bx_in,
      start => VMSMER_D3PHID_start
  );

  LATCH_VMSMER_D3PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D3PHID_bx
  );

  VMSMER_D3PHID : entity work.VMSMER_D3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D3PHID_bx,
      valid        => AS_D3PHIDin_valid,
      index        => AS_D3PHIDin_index,
      allStub_data_V        => AS_D3PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D3PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D3PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D3PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIDn2_din
  );

  VMSMER_D4PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D4PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D4PHIA_bx_in,
      start => VMSMER_D4PHIA_start,
      enb   => AS_D4PHIAin_enb,
      addra => AS_D4PHIAin_V_readaddr,
      din   => AS_D4PHIAin_V_dout,
      dout  => AS_D4PHIAin_V_as,
      valid  => AS_D4PHIAin_valid,
      index  => AS_D4PHIAin_index(6 downto 0),
      nent  => AS_D4PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIA_bx_in,
      start => VMSMER_D4PHIA_start
  );

  LATCH_VMSMER_D4PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIA_bx
  );

  VMSMER_D4PHIA : entity work.VMSMER_D4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D4PHIA_bx,
      valid        => AS_D4PHIAin_valid,
      index        => AS_D4PHIAin_index,
      allStub_data_V        => AS_D4PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D4PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D4PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D4PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIAn2_din
  );

  VMSMER_D4PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D4PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D4PHIB_bx_in,
      start => VMSMER_D4PHIB_start,
      enb   => AS_D4PHIBin_enb,
      addra => AS_D4PHIBin_V_readaddr,
      din   => AS_D4PHIBin_V_dout,
      dout  => AS_D4PHIBin_V_as,
      valid  => AS_D4PHIBin_valid,
      index  => AS_D4PHIBin_index(6 downto 0),
      nent  => AS_D4PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIB_bx_in,
      start => VMSMER_D4PHIB_start
  );

  LATCH_VMSMER_D4PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIB_bx
  );

  VMSMER_D4PHIB : entity work.VMSMER_D4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D4PHIB_bx,
      valid        => AS_D4PHIBin_valid,
      index        => AS_D4PHIBin_index,
      allStub_data_V        => AS_D4PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D4PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D4PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D4PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIBn2_din
  );

  VMSMER_D4PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D4PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D4PHIC_bx_in,
      start => VMSMER_D4PHIC_start,
      enb   => AS_D4PHICin_enb,
      addra => AS_D4PHICin_V_readaddr,
      din   => AS_D4PHICin_V_dout,
      dout  => AS_D4PHICin_V_as,
      valid  => AS_D4PHICin_valid,
      index  => AS_D4PHICin_index(6 downto 0),
      nent  => AS_D4PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIC_bx_in,
      start => VMSMER_D4PHIC_start
  );

  LATCH_VMSMER_D4PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHIC_bx
  );

  VMSMER_D4PHIC : entity work.VMSMER_D4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D4PHIC_bx,
      valid        => AS_D4PHICin_valid,
      index        => AS_D4PHICin_index,
      allStub_data_V        => AS_D4PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D4PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D4PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D4PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHICn2_din
  );

  VMSMER_D4PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D4PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D4PHID_bx_in,
      start => VMSMER_D4PHID_start,
      enb   => AS_D4PHIDin_enb,
      addra => AS_D4PHIDin_V_readaddr,
      din   => AS_D4PHIDin_V_dout,
      dout  => AS_D4PHIDin_V_as,
      valid  => AS_D4PHIDin_valid,
      index  => AS_D4PHIDin_index(6 downto 0),
      nent  => AS_D4PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHID_bx_in,
      start => VMSMER_D4PHID_start
  );

  LATCH_VMSMER_D4PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D4PHID_bx
  );

  VMSMER_D4PHID : entity work.VMSMER_D4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D4PHID_bx,
      valid        => AS_D4PHIDin_valid,
      index        => AS_D4PHIDin_index,
      allStub_data_V        => AS_D4PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D4PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D4PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D4PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIDn2_din
  );

  VMSMER_D5PHIA_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D5PHIA_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D5PHIA_bx_in,
      start => VMSMER_D5PHIA_start,
      enb   => AS_D5PHIAin_enb,
      addra => AS_D5PHIAin_V_readaddr,
      din   => AS_D5PHIAin_V_dout,
      dout  => AS_D5PHIAin_V_as,
      valid  => AS_D5PHIAin_valid,
      index  => AS_D5PHIAin_index(6 downto 0),
      nent  => AS_D5PHIAin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIA_bx_in,
      start => VMSMER_D5PHIA_start
  );

  LATCH_VMSMER_D5PHIA_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIA_bx
  );

  VMSMER_D5PHIA : entity work.VMSMER_D5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D5PHIA_bx,
      valid        => AS_D5PHIAin_valid,
      index        => AS_D5PHIAin_index,
      allStub_data_V        => AS_D5PHIAin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D5PHIAn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D5PHIAn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D5PHIAn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIAn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIAn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIAn2_din
  );

  VMSMER_D5PHIB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D5PHIB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D5PHIB_bx_in,
      start => VMSMER_D5PHIB_start,
      enb   => AS_D5PHIBin_enb,
      addra => AS_D5PHIBin_V_readaddr,
      din   => AS_D5PHIBin_V_dout,
      dout  => AS_D5PHIBin_V_as,
      valid  => AS_D5PHIBin_valid,
      index  => AS_D5PHIBin_index(6 downto 0),
      nent  => AS_D5PHIBin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIB_bx_in,
      start => VMSMER_D5PHIB_start
  );

  LATCH_VMSMER_D5PHIB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIB_bx
  );

  VMSMER_D5PHIB : entity work.VMSMER_D5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D5PHIB_bx,
      valid        => AS_D5PHIBin_valid,
      index        => AS_D5PHIBin_index,
      allStub_data_V        => AS_D5PHIBin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D5PHIBn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D5PHIBn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D5PHIBn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIBn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIBn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIBn2_din
  );

  VMSMER_D5PHIC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D5PHIC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D5PHIC_bx_in,
      start => VMSMER_D5PHIC_start,
      enb   => AS_D5PHICin_enb,
      addra => AS_D5PHICin_V_readaddr,
      din   => AS_D5PHICin_V_dout,
      dout  => AS_D5PHICin_V_as,
      valid  => AS_D5PHICin_valid,
      index  => AS_D5PHICin_index(6 downto 0),
      nent  => AS_D5PHICin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIC_bx_in,
      start => VMSMER_D5PHIC_start
  );

  LATCH_VMSMER_D5PHIC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHIC_bx
  );

  VMSMER_D5PHIC : entity work.VMSMER_D5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D5PHIC_bx,
      valid        => AS_D5PHICin_valid,
      index        => AS_D5PHICin_index,
      allStub_data_V        => AS_D5PHICin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D5PHICn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D5PHICn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D5PHICn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHICn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHICn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHICn2_din
  );

  VMSMER_D5PHID_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 36,
      NAME    => "VMSMER_D5PHID_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => VMSMER_D5PHID_bx_in,
      start => VMSMER_D5PHID_start,
      enb   => AS_D5PHIDin_enb,
      addra => AS_D5PHIDin_V_readaddr,
      din   => AS_D5PHIDin_V_dout,
      dout  => AS_D5PHIDin_V_as,
      valid  => AS_D5PHIDin_valid,
      index  => AS_D5PHIDin_index(6 downto 0),
      nent  => AS_D5PHIDin_AV_dout_nent,
      mask  => (others => (others => '1'))
    );

  LATCH_VMSMER_D5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHID_bx_in,
      start => VMSMER_D5PHID_start
  );

  LATCH_VMSMER_D5PHID_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => VMSMER_D5PHID_bx
  );

  VMSMER_D5PHID : entity work.VMSMER_D5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      bx_V          => VMSMER_D5PHID_bx,
      valid        => AS_D5PHIDin_valid,
      index        => AS_D5PHIDin_index,
      allStub_data_V        => AS_D5PHIDin_V_as,
      memoryME_0_dataarray_0_data_V_ce0       => open,
      memoryME_0_dataarray_0_data_V_we0       => VMSME_D5PHIDn2_wea,
      memoryME_0_dataarray_0_data_V_address0  => VMSME_D5PHIDn2_writeaddr,
      memoryME_0_dataarray_0_data_V_d0        => VMSME_D5PHIDn2_din,
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIDn2_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIDn2_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIDn2_din
  );

  PC_L1L2ABC_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2ABC_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2ABC_bx_in,
      start => PC_L1L2ABC_start,
      enb   => MPAR_L1L2ABCin_enb,
      addra => MPAR_L1L2ABCin_V_readaddr,
      din   => MPAR_L1L2ABCin_V_dout,
      dout  => MPAR_L1L2ABCin_V_tpar,
      valid  => MPAR_L1L2ABCin_valid,
      index  => MPAR_L1L2ABCin_trackletindex,
      nent  => MPAR_L1L2ABCin_AV_dout_nent,
      mask  => MPAR_L1L2ABCin_AV_dout_mask
    );

  LATCH_PC_VMSMER: entity work.tf_pipeline_slr_xing
      generic map (
        NUM_SLR       => 3,
        DELAY         => (2, 119, 2),
        USE_SRL       => (false, true, false)
      )
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_bx_out,
      start => PC_done
  );

  LATCH_PC_L1L2ABC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2ABC_bx_in,
      start => PC_L1L2ABC_start
  );

  LATCH_PC_L1L2ABC_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2ABC_bx
  );

  PC_L1L2ABC : entity work.PC_L1L2ABC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2ABC_bx,
      valid        => MPAR_L1L2ABCin_valid,
      trackletindex_V        => MPAR_L1L2ABCin_trackletindex,
      tpar_data_V        => MPAR_L1L2ABCin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2ABC_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2ABC_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2ABC_din,
      projout_barrel_ps_12_dataarray_data_V_ce0       => open,
      projout_barrel_ps_12_dataarray_data_V_we0       => MPROJ_L1L2ABC_L3PHIA_wea,
      projout_barrel_ps_12_dataarray_data_V_address0  => MPROJ_L1L2ABC_L3PHIA_writeaddr,
      projout_barrel_ps_12_dataarray_data_V_d0        => MPROJ_L1L2ABC_L3PHIA_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L1L2ABC_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L1L2ABC_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L1L2ABC_L3PHIB_din,
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => MPROJ_L1L2ABC_L4PHIA_wea,
      projout_barrel_2s_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L4PHIA_writeaddr,
      projout_barrel_2s_0_dataarray_data_V_d0        => MPROJ_L1L2ABC_L4PHIA_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L1L2ABC_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L1L2ABC_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L1L2ABC_L4PHIB_din,
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => MPROJ_L1L2ABC_L5PHIA_wea,
      projout_barrel_2s_4_dataarray_data_V_address0  => MPROJ_L1L2ABC_L5PHIA_writeaddr,
      projout_barrel_2s_4_dataarray_data_V_d0        => MPROJ_L1L2ABC_L5PHIA_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L1L2ABC_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L1L2ABC_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L1L2ABC_L5PHIB_din,
      projout_barrel_2s_8_dataarray_data_V_ce0       => open,
      projout_barrel_2s_8_dataarray_data_V_we0       => MPROJ_L1L2ABC_L6PHIA_wea,
      projout_barrel_2s_8_dataarray_data_V_address0  => MPROJ_L1L2ABC_L6PHIA_writeaddr,
      projout_barrel_2s_8_dataarray_data_V_d0        => MPROJ_L1L2ABC_L6PHIA_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L1L2ABC_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L1L2ABC_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L1L2ABC_L6PHIB_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_L1L2ABC_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_L1L2ABC_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L1L2ABC_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L1L2ABC_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L1L2ABC_D1PHIB_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L1L2ABC_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L1L2ABC_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L1L2ABC_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1L2ABC_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1L2ABC_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1L2ABC_D2PHIB_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L1L2ABC_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L1L2ABC_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L1L2ABC_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1L2ABC_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1L2ABC_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1L2ABC_D3PHIB_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L1L2ABC_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L1L2ABC_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L1L2ABC_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1L2ABC_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1L2ABC_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1L2ABC_D4PHIB_din
  );

  PC_L1L2DE_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2DE_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2DE_bx_in,
      start => PC_L1L2DE_start,
      enb   => MPAR_L1L2DEin_enb,
      addra => MPAR_L1L2DEin_V_readaddr,
      din   => MPAR_L1L2DEin_V_dout,
      dout  => MPAR_L1L2DEin_V_tpar,
      valid  => MPAR_L1L2DEin_valid,
      index  => MPAR_L1L2DEin_trackletindex,
      nent  => MPAR_L1L2DEin_AV_dout_nent,
      mask  => MPAR_L1L2DEin_AV_dout_mask
    );

  LATCH_PC_L1L2DE: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2DE_bx_in,
      start => PC_L1L2DE_start
  );

  LATCH_PC_L1L2DE_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2DE_bx
  );

  PC_L1L2DE : entity work.PC_L1L2DE
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2DE_bx,
      valid        => MPAR_L1L2DEin_valid,
      trackletindex_V        => MPAR_L1L2DEin_trackletindex,
      tpar_data_V        => MPAR_L1L2DEin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2DE_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2DE_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2DE_din,
      projout_barrel_ps_12_dataarray_data_V_ce0       => open,
      projout_barrel_ps_12_dataarray_data_V_we0       => MPROJ_L1L2DE_L3PHIA_wea,
      projout_barrel_ps_12_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIA_writeaddr,
      projout_barrel_ps_12_dataarray_data_V_d0        => MPROJ_L1L2DE_L3PHIA_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L1L2DE_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L1L2DE_L3PHIB_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L1L2DE_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L1L2DE_L3PHIC_din,
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => MPROJ_L1L2DE_L4PHIA_wea,
      projout_barrel_2s_0_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIA_writeaddr,
      projout_barrel_2s_0_dataarray_data_V_d0        => MPROJ_L1L2DE_L4PHIA_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L1L2DE_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L1L2DE_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L1L2DE_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L1L2DE_L4PHIC_din,
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => MPROJ_L1L2DE_L5PHIA_wea,
      projout_barrel_2s_4_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIA_writeaddr,
      projout_barrel_2s_4_dataarray_data_V_d0        => MPROJ_L1L2DE_L5PHIA_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L1L2DE_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L1L2DE_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L1L2DE_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L1L2DE_L5PHIC_din,
      projout_barrel_2s_8_dataarray_data_V_ce0       => open,
      projout_barrel_2s_8_dataarray_data_V_we0       => MPROJ_L1L2DE_L6PHIA_wea,
      projout_barrel_2s_8_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIA_writeaddr,
      projout_barrel_2s_8_dataarray_data_V_d0        => MPROJ_L1L2DE_L6PHIA_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L1L2DE_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L1L2DE_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L1L2DE_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L1L2DE_L6PHIC_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_L1L2DE_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_L1L2DE_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L1L2DE_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L1L2DE_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L1L2DE_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L1L2DE_D1PHIC_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L1L2DE_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L1L2DE_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1L2DE_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1L2DE_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1L2DE_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1L2DE_D2PHIC_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L1L2DE_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L1L2DE_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1L2DE_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1L2DE_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1L2DE_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1L2DE_D3PHIC_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L1L2DE_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L1L2DE_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1L2DE_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1L2DE_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1L2DE_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1L2DE_D4PHIC_din
  );

  PC_L1L2F_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2F_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2F_bx_in,
      start => PC_L1L2F_start,
      enb   => MPAR_L1L2Fin_enb,
      addra => MPAR_L1L2Fin_V_readaddr,
      din   => MPAR_L1L2Fin_V_dout,
      dout  => MPAR_L1L2Fin_V_tpar,
      valid  => MPAR_L1L2Fin_valid,
      index  => MPAR_L1L2Fin_trackletindex,
      nent  => MPAR_L1L2Fin_AV_dout_nent,
      mask  => MPAR_L1L2Fin_AV_dout_mask
    );

  LATCH_PC_L1L2F: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2F_bx_in,
      start => PC_L1L2F_start
  );

  LATCH_PC_L1L2F_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2F_bx
  );

  PC_L1L2F : entity work.PC_L1L2F
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2F_bx,
      valid        => MPAR_L1L2Fin_valid,
      trackletindex_V        => MPAR_L1L2Fin_trackletindex,
      tpar_data_V        => MPAR_L1L2Fin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2F_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2F_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2F_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L1L2F_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L1L2F_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L1L2F_L3PHIB_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L1L2F_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L1L2F_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L1L2F_L3PHIC_din,
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => MPROJ_L1L2F_L4PHIA_wea,
      projout_barrel_2s_0_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIA_writeaddr,
      projout_barrel_2s_0_dataarray_data_V_d0        => MPROJ_L1L2F_L4PHIA_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L1L2F_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L1L2F_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L1L2F_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L1L2F_L4PHIC_din,
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => MPROJ_L1L2F_L5PHIA_wea,
      projout_barrel_2s_4_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIA_writeaddr,
      projout_barrel_2s_4_dataarray_data_V_d0        => MPROJ_L1L2F_L5PHIA_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L1L2F_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L1L2F_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L1L2F_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L1L2F_L5PHIC_din,
      projout_barrel_2s_8_dataarray_data_V_ce0       => open,
      projout_barrel_2s_8_dataarray_data_V_we0       => MPROJ_L1L2F_L6PHIA_wea,
      projout_barrel_2s_8_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIA_writeaddr,
      projout_barrel_2s_8_dataarray_data_V_d0        => MPROJ_L1L2F_L6PHIA_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L1L2F_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L1L2F_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L1L2F_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L1L2F_L6PHIC_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_L1L2F_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_L1L2F_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L1L2F_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L1L2F_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L1L2F_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L1L2F_D1PHIC_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L1L2F_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L1L2F_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1L2F_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1L2F_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1L2F_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1L2F_D2PHIC_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L1L2F_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L1L2F_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1L2F_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1L2F_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1L2F_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1L2F_D3PHIC_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L1L2F_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L1L2F_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1L2F_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1L2F_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1L2F_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1L2F_D4PHIC_din
  );

  PC_L1L2G_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2G_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2G_bx_in,
      start => PC_L1L2G_start,
      enb   => MPAR_L1L2Gin_enb,
      addra => MPAR_L1L2Gin_V_readaddr,
      din   => MPAR_L1L2Gin_V_dout,
      dout  => MPAR_L1L2Gin_V_tpar,
      valid  => MPAR_L1L2Gin_valid,
      index  => MPAR_L1L2Gin_trackletindex,
      nent  => MPAR_L1L2Gin_AV_dout_nent,
      mask  => MPAR_L1L2Gin_AV_dout_mask
    );

  LATCH_PC_L1L2G: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2G_bx_in,
      start => PC_L1L2G_start
  );

  LATCH_PC_L1L2G_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2G_bx
  );

  PC_L1L2G : entity work.PC_L1L2G
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2G_bx,
      valid        => MPAR_L1L2Gin_valid,
      trackletindex_V        => MPAR_L1L2Gin_trackletindex,
      tpar_data_V        => MPAR_L1L2Gin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2G_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2G_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2G_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L1L2G_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L1L2G_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L1L2G_L3PHIB_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L1L2G_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L1L2G_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L1L2G_L3PHIC_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L1L2G_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L1L2G_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L1L2G_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L1L2G_L4PHIC_din,
      projout_barrel_2s_3_dataarray_data_V_ce0       => open,
      projout_barrel_2s_3_dataarray_data_V_we0       => MPROJ_L1L2G_L4PHID_wea,
      projout_barrel_2s_3_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHID_writeaddr,
      projout_barrel_2s_3_dataarray_data_V_d0        => MPROJ_L1L2G_L4PHID_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L1L2G_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L1L2G_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L1L2G_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L1L2G_L5PHIC_din,
      projout_barrel_2s_7_dataarray_data_V_ce0       => open,
      projout_barrel_2s_7_dataarray_data_V_we0       => MPROJ_L1L2G_L5PHID_wea,
      projout_barrel_2s_7_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHID_writeaddr,
      projout_barrel_2s_7_dataarray_data_V_d0        => MPROJ_L1L2G_L5PHID_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L1L2G_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L1L2G_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L1L2G_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L1L2G_L6PHIC_din,
      projout_barrel_2s_11_dataarray_data_V_ce0       => open,
      projout_barrel_2s_11_dataarray_data_V_we0       => MPROJ_L1L2G_L6PHID_wea,
      projout_barrel_2s_11_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHID_writeaddr,
      projout_barrel_2s_11_dataarray_data_V_d0        => MPROJ_L1L2G_L6PHID_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L1L2G_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L1L2G_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L1L2G_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L1L2G_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_L1L2G_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_L1L2G_D1PHID_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1L2G_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1L2G_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1L2G_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1L2G_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L1L2G_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L1L2G_D2PHID_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1L2G_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1L2G_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1L2G_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1L2G_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L1L2G_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L1L2G_D3PHID_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1L2G_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1L2G_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1L2G_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1L2G_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L1L2G_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L1L2G_D4PHID_din
  );

  PC_L1L2HI_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2HI_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2HI_bx_in,
      start => PC_L1L2HI_start,
      enb   => MPAR_L1L2HIin_enb,
      addra => MPAR_L1L2HIin_V_readaddr,
      din   => MPAR_L1L2HIin_V_dout,
      dout  => MPAR_L1L2HIin_V_tpar,
      valid  => MPAR_L1L2HIin_valid,
      index  => MPAR_L1L2HIin_trackletindex,
      nent  => MPAR_L1L2HIin_AV_dout_nent,
      mask  => MPAR_L1L2HIin_AV_dout_mask
    );

  LATCH_PC_L1L2HI: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2HI_bx_in,
      start => PC_L1L2HI_start
  );

  LATCH_PC_L1L2HI_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2HI_bx
  );

  PC_L1L2HI : entity work.PC_L1L2HI
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2HI_bx,
      valid        => MPAR_L1L2HIin_valid,
      trackletindex_V        => MPAR_L1L2HIin_trackletindex,
      tpar_data_V        => MPAR_L1L2HIin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2HI_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2HI_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2HI_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L1L2HI_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L1L2HI_L3PHIB_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L1L2HI_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L1L2HI_L3PHIC_din,
      projout_barrel_ps_15_dataarray_data_V_ce0       => open,
      projout_barrel_ps_15_dataarray_data_V_we0       => MPROJ_L1L2HI_L3PHID_wea,
      projout_barrel_ps_15_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHID_writeaddr,
      projout_barrel_ps_15_dataarray_data_V_d0        => MPROJ_L1L2HI_L3PHID_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L1L2HI_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L1L2HI_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L1L2HI_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L1L2HI_L4PHIC_din,
      projout_barrel_2s_3_dataarray_data_V_ce0       => open,
      projout_barrel_2s_3_dataarray_data_V_we0       => MPROJ_L1L2HI_L4PHID_wea,
      projout_barrel_2s_3_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHID_writeaddr,
      projout_barrel_2s_3_dataarray_data_V_d0        => MPROJ_L1L2HI_L4PHID_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L1L2HI_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L1L2HI_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L1L2HI_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L1L2HI_L5PHIC_din,
      projout_barrel_2s_7_dataarray_data_V_ce0       => open,
      projout_barrel_2s_7_dataarray_data_V_we0       => MPROJ_L1L2HI_L5PHID_wea,
      projout_barrel_2s_7_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHID_writeaddr,
      projout_barrel_2s_7_dataarray_data_V_d0        => MPROJ_L1L2HI_L5PHID_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L1L2HI_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L1L2HI_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L1L2HI_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L1L2HI_L6PHIC_din,
      projout_barrel_2s_11_dataarray_data_V_ce0       => open,
      projout_barrel_2s_11_dataarray_data_V_we0       => MPROJ_L1L2HI_L6PHID_wea,
      projout_barrel_2s_11_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHID_writeaddr,
      projout_barrel_2s_11_dataarray_data_V_d0        => MPROJ_L1L2HI_L6PHID_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L1L2HI_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L1L2HI_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L1L2HI_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L1L2HI_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_L1L2HI_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_L1L2HI_D1PHID_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1L2HI_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1L2HI_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1L2HI_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1L2HI_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L1L2HI_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L1L2HI_D2PHID_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1L2HI_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1L2HI_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1L2HI_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1L2HI_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L1L2HI_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L1L2HI_D3PHID_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1L2HI_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1L2HI_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1L2HI_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1L2HI_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L1L2HI_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L1L2HI_D4PHID_din
  );

  PC_L1L2JKL_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1L2JKL_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1L2JKL_bx_in,
      start => PC_L1L2JKL_start,
      enb   => MPAR_L1L2JKLin_enb,
      addra => MPAR_L1L2JKLin_V_readaddr,
      din   => MPAR_L1L2JKLin_V_dout,
      dout  => MPAR_L1L2JKLin_V_tpar,
      valid  => MPAR_L1L2JKLin_valid,
      index  => MPAR_L1L2JKLin_trackletindex,
      nent  => MPAR_L1L2JKLin_AV_dout_nent,
      mask  => MPAR_L1L2JKLin_AV_dout_mask
    );

  LATCH_PC_L1L2JKL: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1L2JKL_bx_in,
      start => PC_L1L2JKL_start
  );

  LATCH_PC_L1L2JKL_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1L2JKL_bx
  );

  PC_L1L2JKL : entity work.PC_L1L2JKL
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1L2JKL_bx,
      valid        => MPAR_L1L2JKLin_valid,
      trackletindex_V        => MPAR_L1L2JKLin_trackletindex,
      tpar_data_V        => MPAR_L1L2JKLin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1L2JKL_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1L2JKL_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1L2JKL_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L1L2JKL_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L1L2JKL_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L1L2JKL_L3PHIC_din,
      projout_barrel_ps_15_dataarray_data_V_ce0       => open,
      projout_barrel_ps_15_dataarray_data_V_we0       => MPROJ_L1L2JKL_L3PHID_wea,
      projout_barrel_ps_15_dataarray_data_V_address0  => MPROJ_L1L2JKL_L3PHID_writeaddr,
      projout_barrel_ps_15_dataarray_data_V_d0        => MPROJ_L1L2JKL_L3PHID_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L1L2JKL_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L1L2JKL_L4PHIC_din,
      projout_barrel_2s_3_dataarray_data_V_ce0       => open,
      projout_barrel_2s_3_dataarray_data_V_we0       => MPROJ_L1L2JKL_L4PHID_wea,
      projout_barrel_2s_3_dataarray_data_V_address0  => MPROJ_L1L2JKL_L4PHID_writeaddr,
      projout_barrel_2s_3_dataarray_data_V_d0        => MPROJ_L1L2JKL_L4PHID_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L1L2JKL_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L1L2JKL_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L1L2JKL_L5PHIC_din,
      projout_barrel_2s_7_dataarray_data_V_ce0       => open,
      projout_barrel_2s_7_dataarray_data_V_we0       => MPROJ_L1L2JKL_L5PHID_wea,
      projout_barrel_2s_7_dataarray_data_V_address0  => MPROJ_L1L2JKL_L5PHID_writeaddr,
      projout_barrel_2s_7_dataarray_data_V_d0        => MPROJ_L1L2JKL_L5PHID_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L1L2JKL_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L1L2JKL_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L1L2JKL_L6PHIC_din,
      projout_barrel_2s_11_dataarray_data_V_ce0       => open,
      projout_barrel_2s_11_dataarray_data_V_we0       => MPROJ_L1L2JKL_L6PHID_wea,
      projout_barrel_2s_11_dataarray_data_V_address0  => MPROJ_L1L2JKL_L6PHID_writeaddr,
      projout_barrel_2s_11_dataarray_data_V_d0        => MPROJ_L1L2JKL_L6PHID_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L1L2JKL_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L1L2JKL_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_L1L2JKL_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_L1L2JKL_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_L1L2JKL_D1PHID_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1L2JKL_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1L2JKL_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1L2JKL_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L1L2JKL_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L1L2JKL_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L1L2JKL_D2PHID_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1L2JKL_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1L2JKL_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1L2JKL_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L1L2JKL_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L1L2JKL_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L1L2JKL_D3PHID_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1L2JKL_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1L2JKL_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1L2JKL_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L1L2JKL_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L1L2JKL_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L1L2JKL_D4PHID_din
  );

  PC_L2L3ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L2L3ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L2L3ABCD_bx_in,
      start => PC_L2L3ABCD_start,
      enb   => MPAR_L2L3ABCDin_enb,
      addra => MPAR_L2L3ABCDin_V_readaddr,
      din   => MPAR_L2L3ABCDin_V_dout,
      dout  => MPAR_L2L3ABCDin_V_tpar,
      valid  => MPAR_L2L3ABCDin_valid,
      index  => MPAR_L2L3ABCDin_trackletindex,
      nent  => MPAR_L2L3ABCDin_AV_dout_nent,
      mask  => MPAR_L2L3ABCDin_AV_dout_mask
    );

  LATCH_PC_L2L3ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L2L3ABCD_bx_in,
      start => PC_L2L3ABCD_start
  );

  LATCH_PC_L2L3ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L2L3ABCD_bx
  );

  PC_L2L3ABCD : entity work.PC_L2L3ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L2L3ABCD_bx,
      valid        => MPAR_L2L3ABCDin_valid,
      trackletindex_V        => MPAR_L2L3ABCDin_trackletindex,
      tpar_data_V        => MPAR_L2L3ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L2L3ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_L2L3ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L2L3ABCD_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L1PHIH_din,
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L4PHIA_wea,
      projout_barrel_2s_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIA_writeaddr,
      projout_barrel_2s_0_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L4PHIA_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L4PHIC_din,
      projout_barrel_2s_3_dataarray_data_V_ce0       => open,
      projout_barrel_2s_3_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L4PHID_wea,
      projout_barrel_2s_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHID_writeaddr,
      projout_barrel_2s_3_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L4PHID_din,
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L5PHIA_wea,
      projout_barrel_2s_4_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIA_writeaddr,
      projout_barrel_2s_4_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L5PHIA_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L5PHIC_din,
      projout_barrel_2s_7_dataarray_data_V_ce0       => open,
      projout_barrel_2s_7_dataarray_data_V_we0       => MPROJ_L2L3ABCD_L5PHID_wea,
      projout_barrel_2s_7_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHID_writeaddr,
      projout_barrel_2s_7_dataarray_data_V_d0        => MPROJ_L2L3ABCD_L5PHID_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D1PHID_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D2PHID_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D3PHID_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L2L3ABCD_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L2L3ABCD_D4PHID_din
  );

  PC_L3L4AB_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L3L4AB_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L3L4AB_bx_in,
      start => PC_L3L4AB_start,
      enb   => MPAR_L3L4ABin_enb,
      addra => MPAR_L3L4ABin_V_readaddr,
      din   => MPAR_L3L4ABin_V_dout,
      dout  => MPAR_L3L4ABin_V_tpar,
      valid  => MPAR_L3L4ABin_valid,
      index  => MPAR_L3L4ABin_trackletindex,
      nent  => MPAR_L3L4ABin_AV_dout_nent,
      mask  => MPAR_L3L4ABin_AV_dout_mask
    );

  LATCH_PC_L3L4AB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L3L4AB_bx_in,
      start => PC_L3L4AB_start
  );

  LATCH_PC_L3L4AB_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L3L4AB_bx
  );

  PC_L3L4AB : entity work.PC_L3L4AB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L3L4AB_bx,
      valid        => MPAR_L3L4ABin_valid,
      trackletindex_V        => MPAR_L3L4ABin_trackletindex,
      tpar_data_V        => MPAR_L3L4ABin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L3L4AB_wea,
      tparout_dataarray_data_V_address0  => MPAR_L3L4AB_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L3L4AB_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_L3L4AB_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_L3L4AB_L1PHIF_din,
      projout_barrel_ps_8_dataarray_data_V_ce0       => open,
      projout_barrel_ps_8_dataarray_data_V_we0       => MPROJ_L3L4AB_L2PHIA_wea,
      projout_barrel_ps_8_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIA_writeaddr,
      projout_barrel_ps_8_dataarray_data_V_d0        => MPROJ_L3L4AB_L2PHIA_din,
      projout_barrel_ps_9_dataarray_data_V_ce0       => open,
      projout_barrel_ps_9_dataarray_data_V_we0       => MPROJ_L3L4AB_L2PHIB_wea,
      projout_barrel_ps_9_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIB_writeaddr,
      projout_barrel_ps_9_dataarray_data_V_d0        => MPROJ_L3L4AB_L2PHIB_din,
      projout_barrel_ps_10_dataarray_data_V_ce0       => open,
      projout_barrel_ps_10_dataarray_data_V_we0       => MPROJ_L3L4AB_L2PHIC_wea,
      projout_barrel_ps_10_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIC_writeaddr,
      projout_barrel_ps_10_dataarray_data_V_d0        => MPROJ_L3L4AB_L2PHIC_din,
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => MPROJ_L3L4AB_L5PHIA_wea,
      projout_barrel_2s_4_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIA_writeaddr,
      projout_barrel_2s_4_dataarray_data_V_d0        => MPROJ_L3L4AB_L5PHIA_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L3L4AB_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L3L4AB_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L3L4AB_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L3L4AB_L5PHIC_din,
      projout_barrel_2s_8_dataarray_data_V_ce0       => open,
      projout_barrel_2s_8_dataarray_data_V_we0       => MPROJ_L3L4AB_L6PHIA_wea,
      projout_barrel_2s_8_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIA_writeaddr,
      projout_barrel_2s_8_dataarray_data_V_d0        => MPROJ_L3L4AB_L6PHIA_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L3L4AB_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L3L4AB_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L3L4AB_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L3L4AB_L6PHIC_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_L3L4AB_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_L3L4AB_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L3L4AB_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L3L4AB_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L3L4AB_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L3L4AB_D1PHIC_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L3L4AB_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L3L4AB_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L3L4AB_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L3L4AB_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L3L4AB_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L3L4AB_D2PHIC_din
  );

  PC_L3L4CD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L3L4CD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L3L4CD_bx_in,
      start => PC_L3L4CD_start,
      enb   => MPAR_L3L4CDin_enb,
      addra => MPAR_L3L4CDin_V_readaddr,
      din   => MPAR_L3L4CDin_V_dout,
      dout  => MPAR_L3L4CDin_V_tpar,
      valid  => MPAR_L3L4CDin_valid,
      index  => MPAR_L3L4CDin_trackletindex,
      nent  => MPAR_L3L4CDin_AV_dout_nent,
      mask  => MPAR_L3L4CDin_AV_dout_mask
    );

  LATCH_PC_L3L4CD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L3L4CD_bx_in,
      start => PC_L3L4CD_start
  );

  LATCH_PC_L3L4CD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L3L4CD_bx
  );

  PC_L3L4CD : entity work.PC_L3L4CD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L3L4CD_bx,
      valid        => MPAR_L3L4CDin_valid,
      trackletindex_V        => MPAR_L3L4CDin_trackletindex,
      tpar_data_V        => MPAR_L3L4CDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L3L4CD_wea,
      tparout_dataarray_data_V_address0  => MPAR_L3L4CD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L3L4CD_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_L3L4CD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_L3L4CD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_L3L4CD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_L3L4CD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_L3L4CD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_L3L4CD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_L3L4CD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_L3L4CD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_L3L4CD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_L3L4CD_L1PHIH_din,
      projout_barrel_ps_9_dataarray_data_V_ce0       => open,
      projout_barrel_ps_9_dataarray_data_V_we0       => MPROJ_L3L4CD_L2PHIB_wea,
      projout_barrel_ps_9_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHIB_writeaddr,
      projout_barrel_ps_9_dataarray_data_V_d0        => MPROJ_L3L4CD_L2PHIB_din,
      projout_barrel_ps_10_dataarray_data_V_ce0       => open,
      projout_barrel_ps_10_dataarray_data_V_we0       => MPROJ_L3L4CD_L2PHIC_wea,
      projout_barrel_ps_10_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHIC_writeaddr,
      projout_barrel_ps_10_dataarray_data_V_d0        => MPROJ_L3L4CD_L2PHIC_din,
      projout_barrel_ps_11_dataarray_data_V_ce0       => open,
      projout_barrel_ps_11_dataarray_data_V_we0       => MPROJ_L3L4CD_L2PHID_wea,
      projout_barrel_ps_11_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHID_writeaddr,
      projout_barrel_ps_11_dataarray_data_V_d0        => MPROJ_L3L4CD_L2PHID_din,
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => MPROJ_L3L4CD_L5PHIB_wea,
      projout_barrel_2s_5_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHIB_writeaddr,
      projout_barrel_2s_5_dataarray_data_V_d0        => MPROJ_L3L4CD_L5PHIB_din,
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => MPROJ_L3L4CD_L5PHIC_wea,
      projout_barrel_2s_6_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHIC_writeaddr,
      projout_barrel_2s_6_dataarray_data_V_d0        => MPROJ_L3L4CD_L5PHIC_din,
      projout_barrel_2s_7_dataarray_data_V_ce0       => open,
      projout_barrel_2s_7_dataarray_data_V_we0       => MPROJ_L3L4CD_L5PHID_wea,
      projout_barrel_2s_7_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHID_writeaddr,
      projout_barrel_2s_7_dataarray_data_V_d0        => MPROJ_L3L4CD_L5PHID_din,
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => MPROJ_L3L4CD_L6PHIB_wea,
      projout_barrel_2s_9_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHIB_writeaddr,
      projout_barrel_2s_9_dataarray_data_V_d0        => MPROJ_L3L4CD_L6PHIB_din,
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => MPROJ_L3L4CD_L6PHIC_wea,
      projout_barrel_2s_10_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHIC_writeaddr,
      projout_barrel_2s_10_dataarray_data_V_d0        => MPROJ_L3L4CD_L6PHIC_din,
      projout_barrel_2s_11_dataarray_data_V_ce0       => open,
      projout_barrel_2s_11_dataarray_data_V_we0       => MPROJ_L3L4CD_L6PHID_wea,
      projout_barrel_2s_11_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHID_writeaddr,
      projout_barrel_2s_11_dataarray_data_V_d0        => MPROJ_L3L4CD_L6PHID_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_L3L4CD_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_L3L4CD_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_L3L4CD_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_L3L4CD_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_L3L4CD_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_L3L4CD_D1PHID_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L3L4CD_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L3L4CD_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L3L4CD_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L3L4CD_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L3L4CD_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L3L4CD_D2PHID_din
  );

  PC_L5L6ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L5L6ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L5L6ABCD_bx_in,
      start => PC_L5L6ABCD_start,
      enb   => MPAR_L5L6ABCDin_enb,
      addra => MPAR_L5L6ABCDin_V_readaddr,
      din   => MPAR_L5L6ABCDin_V_dout,
      dout  => MPAR_L5L6ABCDin_V_tpar,
      valid  => MPAR_L5L6ABCDin_valid,
      index  => MPAR_L5L6ABCDin_trackletindex,
      nent  => MPAR_L5L6ABCDin_AV_dout_nent,
      mask  => MPAR_L5L6ABCDin_AV_dout_mask
    );

  LATCH_PC_L5L6ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L5L6ABCD_bx_in,
      start => PC_L5L6ABCD_start
  );

  LATCH_PC_L5L6ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L5L6ABCD_bx
  );

  PC_L5L6ABCD : entity work.PC_L5L6ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L5L6ABCD_bx,
      valid        => MPAR_L5L6ABCDin_valid,
      trackletindex_V        => MPAR_L5L6ABCDin_trackletindex,
      tpar_data_V        => MPAR_L5L6ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L5L6ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_L5L6ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L5L6ABCD_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L1PHIH_din,
      projout_barrel_ps_8_dataarray_data_V_ce0       => open,
      projout_barrel_ps_8_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L2PHIA_wea,
      projout_barrel_ps_8_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIA_writeaddr,
      projout_barrel_ps_8_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L2PHIA_din,
      projout_barrel_ps_9_dataarray_data_V_ce0       => open,
      projout_barrel_ps_9_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L2PHIB_wea,
      projout_barrel_ps_9_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIB_writeaddr,
      projout_barrel_ps_9_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L2PHIB_din,
      projout_barrel_ps_10_dataarray_data_V_ce0       => open,
      projout_barrel_ps_10_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L2PHIC_wea,
      projout_barrel_ps_10_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIC_writeaddr,
      projout_barrel_ps_10_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L2PHIC_din,
      projout_barrel_ps_11_dataarray_data_V_ce0       => open,
      projout_barrel_ps_11_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L2PHID_wea,
      projout_barrel_ps_11_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHID_writeaddr,
      projout_barrel_ps_11_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L2PHID_din,
      projout_barrel_ps_12_dataarray_data_V_ce0       => open,
      projout_barrel_ps_12_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L3PHIA_wea,
      projout_barrel_ps_12_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIA_writeaddr,
      projout_barrel_ps_12_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L3PHIA_din,
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L3PHIB_wea,
      projout_barrel_ps_13_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIB_writeaddr,
      projout_barrel_ps_13_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L3PHIB_din,
      projout_barrel_ps_14_dataarray_data_V_ce0       => open,
      projout_barrel_ps_14_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L3PHIC_wea,
      projout_barrel_ps_14_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIC_writeaddr,
      projout_barrel_ps_14_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L3PHIC_din,
      projout_barrel_ps_15_dataarray_data_V_ce0       => open,
      projout_barrel_ps_15_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L3PHID_wea,
      projout_barrel_ps_15_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHID_writeaddr,
      projout_barrel_ps_15_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L3PHID_din,
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L4PHIA_wea,
      projout_barrel_2s_0_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIA_writeaddr,
      projout_barrel_2s_0_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L4PHIA_din,
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L4PHIB_wea,
      projout_barrel_2s_1_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIB_writeaddr,
      projout_barrel_2s_1_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L4PHIB_din,
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L4PHIC_wea,
      projout_barrel_2s_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIC_writeaddr,
      projout_barrel_2s_2_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L4PHIC_din,
      projout_barrel_2s_3_dataarray_data_V_ce0       => open,
      projout_barrel_2s_3_dataarray_data_V_we0       => MPROJ_L5L6ABCD_L4PHID_wea,
      projout_barrel_2s_3_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHID_writeaddr,
      projout_barrel_2s_3_dataarray_data_V_d0        => MPROJ_L5L6ABCD_L4PHID_din
  );

  PC_D1D2ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_D1D2ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_D1D2ABCD_bx_in,
      start => PC_D1D2ABCD_start,
      enb   => MPAR_D1D2ABCDin_enb,
      addra => MPAR_D1D2ABCDin_V_readaddr,
      din   => MPAR_D1D2ABCDin_V_dout,
      dout  => MPAR_D1D2ABCDin_V_tpar,
      valid  => MPAR_D1D2ABCDin_valid,
      index  => MPAR_D1D2ABCDin_trackletindex,
      nent  => MPAR_D1D2ABCDin_AV_dout_nent,
      mask  => MPAR_D1D2ABCDin_AV_dout_mask
    );

  LATCH_PC_D1D2ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_D1D2ABCD_bx_in,
      start => PC_D1D2ABCD_start
  );

  LATCH_PC_D1D2ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_D1D2ABCD_bx
  );

  PC_D1D2ABCD : entity work.PC_D1D2ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_D1D2ABCD_bx,
      valid        => MPAR_D1D2ABCDin_valid,
      trackletindex_V        => MPAR_D1D2ABCDin_trackletindex,
      tpar_data_V        => MPAR_D1D2ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_D1D2ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_D1D2ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_D1D2ABCD_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L1PHIH_din,
      projout_barrel_ps_8_dataarray_data_V_ce0       => open,
      projout_barrel_ps_8_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L2PHIA_wea,
      projout_barrel_ps_8_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIA_writeaddr,
      projout_barrel_ps_8_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L2PHIA_din,
      projout_barrel_ps_9_dataarray_data_V_ce0       => open,
      projout_barrel_ps_9_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L2PHIB_wea,
      projout_barrel_ps_9_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIB_writeaddr,
      projout_barrel_ps_9_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L2PHIB_din,
      projout_barrel_ps_10_dataarray_data_V_ce0       => open,
      projout_barrel_ps_10_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L2PHIC_wea,
      projout_barrel_ps_10_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIC_writeaddr,
      projout_barrel_ps_10_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L2PHIC_din,
      projout_barrel_ps_11_dataarray_data_V_ce0       => open,
      projout_barrel_ps_11_dataarray_data_V_we0       => MPROJ_D1D2ABCD_L2PHID_wea,
      projout_barrel_ps_11_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHID_writeaddr,
      projout_barrel_ps_11_dataarray_data_V_d0        => MPROJ_D1D2ABCD_L2PHID_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D3PHID_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D4PHID_din,
      projout_disk_16_dataarray_data_V_ce0       => open,
      projout_disk_16_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D5PHIA_wea,
      projout_disk_16_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIA_writeaddr,
      projout_disk_16_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D5PHIA_din,
      projout_disk_17_dataarray_data_V_ce0       => open,
      projout_disk_17_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D5PHIB_wea,
      projout_disk_17_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIB_writeaddr,
      projout_disk_17_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D5PHIB_din,
      projout_disk_18_dataarray_data_V_ce0       => open,
      projout_disk_18_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D5PHIC_wea,
      projout_disk_18_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIC_writeaddr,
      projout_disk_18_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D5PHIC_din,
      projout_disk_19_dataarray_data_V_ce0       => open,
      projout_disk_19_dataarray_data_V_we0       => MPROJ_D1D2ABCD_D5PHID_wea,
      projout_disk_19_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHID_writeaddr,
      projout_disk_19_dataarray_data_V_d0        => MPROJ_D1D2ABCD_D5PHID_din
  );

  PC_D3D4ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_D3D4ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_D3D4ABCD_bx_in,
      start => PC_D3D4ABCD_start,
      enb   => MPAR_D3D4ABCDin_enb,
      addra => MPAR_D3D4ABCDin_V_readaddr,
      din   => MPAR_D3D4ABCDin_V_dout,
      dout  => MPAR_D3D4ABCDin_V_tpar,
      valid  => MPAR_D3D4ABCDin_valid,
      index  => MPAR_D3D4ABCDin_trackletindex,
      nent  => MPAR_D3D4ABCDin_AV_dout_nent,
      mask  => MPAR_D3D4ABCDin_AV_dout_mask
    );

  LATCH_PC_D3D4ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_D3D4ABCD_bx_in,
      start => PC_D3D4ABCD_start
  );

  LATCH_PC_D3D4ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_D3D4ABCD_bx
  );

  PC_D3D4ABCD : entity work.PC_D3D4ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_D3D4ABCD_bx,
      valid        => MPAR_D3D4ABCDin_valid,
      trackletindex_V        => MPAR_D3D4ABCDin_trackletindex,
      tpar_data_V        => MPAR_D3D4ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_D3D4ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_D3D4ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_D3D4ABCD_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_D3D4ABCD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_D3D4ABCD_L1PHIH_din,
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D1PHIA_wea,
      projout_disk_0_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIA_writeaddr,
      projout_disk_0_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D1PHIA_din,
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D1PHIB_wea,
      projout_disk_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIB_writeaddr,
      projout_disk_1_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D1PHIB_din,
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D1PHIC_wea,
      projout_disk_2_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIC_writeaddr,
      projout_disk_2_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D1PHIC_din,
      projout_disk_3_dataarray_data_V_ce0       => open,
      projout_disk_3_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D1PHID_wea,
      projout_disk_3_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHID_writeaddr,
      projout_disk_3_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D1PHID_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D2PHID_din,
      projout_disk_16_dataarray_data_V_ce0       => open,
      projout_disk_16_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D5PHIA_wea,
      projout_disk_16_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIA_writeaddr,
      projout_disk_16_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D5PHIA_din,
      projout_disk_17_dataarray_data_V_ce0       => open,
      projout_disk_17_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D5PHIB_wea,
      projout_disk_17_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIB_writeaddr,
      projout_disk_17_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D5PHIB_din,
      projout_disk_18_dataarray_data_V_ce0       => open,
      projout_disk_18_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D5PHIC_wea,
      projout_disk_18_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIC_writeaddr,
      projout_disk_18_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D5PHIC_din,
      projout_disk_19_dataarray_data_V_ce0       => open,
      projout_disk_19_dataarray_data_V_we0       => MPROJ_D3D4ABCD_D5PHID_wea,
      projout_disk_19_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHID_writeaddr,
      projout_disk_19_dataarray_data_V_d0        => MPROJ_D3D4ABCD_D5PHID_din
  );

  PC_L1D1ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1D1ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1D1ABCD_bx_in,
      start => PC_L1D1ABCD_start,
      enb   => MPAR_L1D1ABCDin_enb,
      addra => MPAR_L1D1ABCDin_V_readaddr,
      din   => MPAR_L1D1ABCDin_V_dout,
      dout  => MPAR_L1D1ABCDin_V_tpar,
      valid  => MPAR_L1D1ABCDin_valid,
      index  => MPAR_L1D1ABCDin_trackletindex,
      nent  => MPAR_L1D1ABCDin_AV_dout_nent,
      mask  => MPAR_L1D1ABCDin_AV_dout_mask
    );

  LATCH_PC_L1D1ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1D1ABCD_bx_in,
      start => PC_L1D1ABCD_start
  );

  LATCH_PC_L1D1ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1D1ABCD_bx
  );

  PC_L1D1ABCD : entity work.PC_L1D1ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1D1ABCD_bx,
      valid        => MPAR_L1D1ABCDin_valid,
      trackletindex_V        => MPAR_L1D1ABCDin_trackletindex,
      tpar_data_V        => MPAR_L1D1ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1D1ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1D1ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1D1ABCD_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D2PHIC_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D3PHIC_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D4PHIC_din,
      projout_disk_16_dataarray_data_V_ce0       => open,
      projout_disk_16_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D5PHIA_wea,
      projout_disk_16_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIA_writeaddr,
      projout_disk_16_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D5PHIA_din,
      projout_disk_17_dataarray_data_V_ce0       => open,
      projout_disk_17_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D5PHIB_wea,
      projout_disk_17_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIB_writeaddr,
      projout_disk_17_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D5PHIB_din,
      projout_disk_18_dataarray_data_V_ce0       => open,
      projout_disk_18_dataarray_data_V_we0       => MPROJ_L1D1ABCD_D5PHIC_wea,
      projout_disk_18_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIC_writeaddr,
      projout_disk_18_dataarray_data_V_d0        => MPROJ_L1D1ABCD_D5PHIC_din
  );

  PC_L1D1EFGH_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L1D1EFGH_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L1D1EFGH_bx_in,
      start => PC_L1D1EFGH_start,
      enb   => MPAR_L1D1EFGHin_enb,
      addra => MPAR_L1D1EFGHin_V_readaddr,
      din   => MPAR_L1D1EFGHin_V_dout,
      dout  => MPAR_L1D1EFGHin_V_tpar,
      valid  => MPAR_L1D1EFGHin_valid,
      index  => MPAR_L1D1EFGHin_trackletindex,
      nent  => MPAR_L1D1EFGHin_AV_dout_nent,
      mask  => MPAR_L1D1EFGHin_AV_dout_mask
    );

  LATCH_PC_L1D1EFGH: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L1D1EFGH_bx_in,
      start => PC_L1D1EFGH_start
  );

  LATCH_PC_L1D1EFGH_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L1D1EFGH_bx
  );

  PC_L1D1EFGH : entity work.PC_L1D1EFGH
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L1D1EFGH_bx,
      valid        => MPAR_L1D1EFGHin_valid,
      trackletindex_V        => MPAR_L1D1EFGHin_trackletindex,
      tpar_data_V        => MPAR_L1D1EFGHin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L1D1EFGH_wea,
      tparout_dataarray_data_V_address0  => MPAR_L1D1EFGH_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L1D1EFGH_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D2PHID_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D3PHID_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D4PHID_din,
      projout_disk_17_dataarray_data_V_ce0       => open,
      projout_disk_17_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D5PHIB_wea,
      projout_disk_17_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHIB_writeaddr,
      projout_disk_17_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D5PHIB_din,
      projout_disk_18_dataarray_data_V_ce0       => open,
      projout_disk_18_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D5PHIC_wea,
      projout_disk_18_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHIC_writeaddr,
      projout_disk_18_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D5PHIC_din,
      projout_disk_19_dataarray_data_V_ce0       => open,
      projout_disk_19_dataarray_data_V_we0       => MPROJ_L1D1EFGH_D5PHID_wea,
      projout_disk_19_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHID_writeaddr,
      projout_disk_19_dataarray_data_V_d0        => MPROJ_L1D1EFGH_D5PHID_din
  );

  PC_L2D1ABCD_mem_reader : entity work.mem_reader
    generic map (
      RAM_WIDTH    => 73,
      NUM_TPAGES    => 4,
      NAME    => "PC_L2D1ABCD_mem_reader"
    )
    port map (
      clk    => clk,
      bx    => PC_L2D1ABCD_bx_in,
      start => PC_L2D1ABCD_start,
      enb   => MPAR_L2D1ABCDin_enb,
      addra => MPAR_L2D1ABCDin_V_readaddr,
      din   => MPAR_L2D1ABCDin_V_dout,
      dout  => MPAR_L2D1ABCDin_V_tpar,
      valid  => MPAR_L2D1ABCDin_valid,
      index  => MPAR_L2D1ABCDin_trackletindex,
      nent  => MPAR_L2D1ABCDin_AV_dout_nent,
      mask  => MPAR_L2D1ABCDin_AV_dout_mask
    );

  LATCH_PC_L2D1ABCD: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_start,
      bx_out => PC_bx_in,
      bx => PC_L2D1ABCD_bx_in,
      start => PC_L2D1ABCD_start
  );

  LATCH_PC_L2D1ABCD_BX_GEN: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      bx_out => PC_bx_in,
      bx => PC_L2D1ABCD_bx
  );

  PC_L2D1ABCD : entity work.PC_L2D1ABCD
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => '1',
      bx_V          => PC_L2D1ABCD_bx,
      valid        => MPAR_L2D1ABCDin_valid,
      trackletindex_V        => MPAR_L2D1ABCDin_trackletindex,
      tpar_data_V        => MPAR_L2D1ABCDin_V_tpar,
      tparout_dataarray_data_V_ce0       => open,
      tparout_dataarray_data_V_we0       => MPAR_L2D1ABCD_wea,
      tparout_dataarray_data_V_address0  => MPAR_L2D1ABCD_writeaddr,
      tparout_dataarray_data_V_d0        => MPAR_L2D1ABCD_din,
      projout_barrel_ps_0_dataarray_data_V_ce0       => open,
      projout_barrel_ps_0_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIA_wea,
      projout_barrel_ps_0_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIA_writeaddr,
      projout_barrel_ps_0_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIA_din,
      projout_barrel_ps_1_dataarray_data_V_ce0       => open,
      projout_barrel_ps_1_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIB_wea,
      projout_barrel_ps_1_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIB_writeaddr,
      projout_barrel_ps_1_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIB_din,
      projout_barrel_ps_2_dataarray_data_V_ce0       => open,
      projout_barrel_ps_2_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIC_wea,
      projout_barrel_ps_2_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIC_writeaddr,
      projout_barrel_ps_2_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIC_din,
      projout_barrel_ps_3_dataarray_data_V_ce0       => open,
      projout_barrel_ps_3_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHID_wea,
      projout_barrel_ps_3_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHID_writeaddr,
      projout_barrel_ps_3_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHID_din,
      projout_barrel_ps_4_dataarray_data_V_ce0       => open,
      projout_barrel_ps_4_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIE_wea,
      projout_barrel_ps_4_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIE_writeaddr,
      projout_barrel_ps_4_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIE_din,
      projout_barrel_ps_5_dataarray_data_V_ce0       => open,
      projout_barrel_ps_5_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIF_wea,
      projout_barrel_ps_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIF_writeaddr,
      projout_barrel_ps_5_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIF_din,
      projout_barrel_ps_6_dataarray_data_V_ce0       => open,
      projout_barrel_ps_6_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIG_wea,
      projout_barrel_ps_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIG_writeaddr,
      projout_barrel_ps_6_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIG_din,
      projout_barrel_ps_7_dataarray_data_V_ce0       => open,
      projout_barrel_ps_7_dataarray_data_V_we0       => MPROJ_L2D1ABCD_L1PHIH_wea,
      projout_barrel_ps_7_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIH_writeaddr,
      projout_barrel_ps_7_dataarray_data_V_d0        => MPROJ_L2D1ABCD_L1PHIH_din,
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D2PHIA_wea,
      projout_disk_4_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIA_writeaddr,
      projout_disk_4_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D2PHIA_din,
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D2PHIB_wea,
      projout_disk_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIB_writeaddr,
      projout_disk_5_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D2PHIB_din,
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D2PHIC_wea,
      projout_disk_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIC_writeaddr,
      projout_disk_6_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D2PHIC_din,
      projout_disk_7_dataarray_data_V_ce0       => open,
      projout_disk_7_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D2PHID_wea,
      projout_disk_7_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHID_writeaddr,
      projout_disk_7_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D2PHID_din,
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D3PHIA_wea,
      projout_disk_8_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIA_writeaddr,
      projout_disk_8_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D3PHIA_din,
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D3PHIB_wea,
      projout_disk_9_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIB_writeaddr,
      projout_disk_9_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D3PHIB_din,
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D3PHIC_wea,
      projout_disk_10_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIC_writeaddr,
      projout_disk_10_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D3PHIC_din,
      projout_disk_11_dataarray_data_V_ce0       => open,
      projout_disk_11_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D3PHID_wea,
      projout_disk_11_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHID_writeaddr,
      projout_disk_11_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D3PHID_din,
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D4PHIA_wea,
      projout_disk_12_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIA_writeaddr,
      projout_disk_12_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D4PHIA_din,
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D4PHIB_wea,
      projout_disk_13_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIB_writeaddr,
      projout_disk_13_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D4PHIB_din,
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D4PHIC_wea,
      projout_disk_14_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIC_writeaddr,
      projout_disk_14_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D4PHIC_din,
      projout_disk_15_dataarray_data_V_ce0       => open,
      projout_disk_15_dataarray_data_V_we0       => MPROJ_L2D1ABCD_D4PHID_wea,
      projout_disk_15_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHID_writeaddr,
      projout_disk_15_dataarray_data_V_d0        => MPROJ_L2D1ABCD_D4PHID_din
  );

  LATCH_MP_L1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIA_bx,
      start => MP_L1PHIA_start
  );

  MP_L1PHIA : entity work.MP_L1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => MP_done,
      bx_V          => MP_L1PHIA_bx,
      bx_o_V        => MP_bx_out,
      bx_o_V_ap_vld => open,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIA_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIA_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIA_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIA_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIA_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIA_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIA_din
  );

  LATCH_MP_L1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIB_bx,
      start => MP_L1PHIB_start
  );

  MP_L1PHIB : entity work.MP_L1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIB_din
  );

  LATCH_MP_L1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIC_bx,
      start => MP_L1PHIC_start
  );

  MP_L1PHIC : entity work.MP_L1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIC_din
  );

  LATCH_MP_L1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHID_bx,
      start => MP_L1PHID_start
  );

  MP_L1PHID : entity work.MP_L1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L3L4CD_L1PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L3L4CD_L1PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L3L4CD_L1PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L3L4CD_L1PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L3L4CD_L1PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L5L6ABCD_L1PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L5L6ABCD_L1PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L5L6ABCD_L1PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_L1PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_L1PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_L1PHID_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHID_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHID_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHID_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_L1PHID_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_L1PHID_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_L1PHID_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHID_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHID_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHID_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_L1PHID_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_L1PHID_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_L1PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHID_din
  );

  LATCH_MP_L1PHIE: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIE_bx,
      start => MP_L1PHIE_start
  );

  MP_L1PHIE : entity work.MP_L1PHIE
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIE_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIE_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIE_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIE_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIE_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIE_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIE_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHIE_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIE_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHIE_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHIE_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHIE_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHIE_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L3L4CD_L1PHIE_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIE_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L3L4CD_L1PHIE_V_dout,
      projin_2_mask_0_V                   => MPROJ_L3L4CD_L1PHIE_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L3L4CD_L1PHIE_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L3L4CD_L1PHIE_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIE_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIE_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIE_V_dout,
      projin_3_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIE_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIE_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIE_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIE_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIE_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIE_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIE_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIE_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIE_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIE_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIE_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIE_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIE_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIE_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIE_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIE_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIE_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIE_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIE_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIE_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIE_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIEn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIEn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIEn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIEn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIEn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIEn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIEn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIEn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIEn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIEn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIEn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIEn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIEn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIEn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIEn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIEn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIEn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIEn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIEn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIEn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIEn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIEn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIEn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIEn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIE_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIE_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIE_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIE_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIE_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIE_din
  );

  LATCH_MP_L1PHIF: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIF_bx,
      start => MP_L1PHIF_start
  );

  MP_L1PHIF : entity work.MP_L1PHIF
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIF_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIF_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIF_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIF_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIF_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIF_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIF_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIF_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4AB_L1PHIF_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4AB_L1PHIF_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4AB_L1PHIF_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4AB_L1PHIF_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4AB_L1PHIF_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4AB_L1PHIF_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L3L4CD_L1PHIF_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIF_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L3L4CD_L1PHIF_V_dout,
      projin_2_mask_0_V                   => MPROJ_L3L4CD_L1PHIF_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L3L4CD_L1PHIF_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L3L4CD_L1PHIF_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIF_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIF_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIF_V_dout,
      projin_3_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIF_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIF_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIF_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIF_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIF_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIF_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIF_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIF_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIF_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIF_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIF_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIF_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIF_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIF_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIF_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIF_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIF_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIF_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIF_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIF_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIF_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIFn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIFn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIFn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIFn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIFn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIFn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIFn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIFn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIFn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIFn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIFn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIFn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIFn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIFn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIFn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIFn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIFn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIFn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIFn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIFn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIFn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIFn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIFn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIFn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIF_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIF_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIF_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIF_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIF_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIF_din
  );

  LATCH_MP_L1PHIG: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIG_bx,
      start => MP_L1PHIG_start
  );

  MP_L1PHIG : entity work.MP_L1PHIG
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIG_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIG_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIG_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIG_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIG_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIG_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIG_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIG_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4CD_L1PHIG_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIG_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4CD_L1PHIG_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4CD_L1PHIG_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4CD_L1PHIG_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4CD_L1PHIG_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIG_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIG_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIG_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIG_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIG_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIG_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIG_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIG_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIG_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIG_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIG_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIG_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIG_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIG_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIG_V_dout,
      projin_4_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIG_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIG_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIG_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIG_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIG_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIG_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIG_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIG_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIG_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIGn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIGn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIGn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIGn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIGn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIGn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIGn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIGn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIGn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIGn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIGn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIGn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIGn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIGn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIGn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIGn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIGn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIGn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIGn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIGn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIGn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIGn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIGn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIGn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIG_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIG_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIG_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIG_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIG_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIG_din
  );

  LATCH_MP_L1PHIH: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L1PHIH_bx,
      start => MP_L1PHIH_start
  );

  MP_L1PHIH : entity work.MP_L1PHIH
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L1PHIH_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L1PHIH_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L1PHIH_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L1PHIH_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L1PHIH_V_dout,
      projin_0_mask_0_V                   => MPROJ_L2L3ABCD_L1PHIH_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L2L3ABCD_L1PHIH_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L2L3ABCD_L1PHIH_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4CD_L1PHIH_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4CD_L1PHIH_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4CD_L1PHIH_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4CD_L1PHIH_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4CD_L1PHIH_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4CD_L1PHIH_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L1PHIH_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L1PHIH_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L1PHIH_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L1PHIH_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L1PHIH_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L1PHIH_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L1PHIH_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L1PHIH_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L1PHIH_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L1PHIH_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L1PHIH_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L1PHIH_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_L1PHIH_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D3D4ABCD_L1PHIH_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D3D4ABCD_L1PHIH_V_dout,
      projin_4_mask_0_V                   => MPROJ_D3D4ABCD_L1PHIH_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D3D4ABCD_L1PHIH_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D3D4ABCD_L1PHIH_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_L1PHIH_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2D1ABCD_L1PHIH_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2D1ABCD_L1PHIH_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2D1ABCD_L1PHIH_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2D1ABCD_L1PHIH_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2D1ABCD_L1PHIH_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L1PHIHn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L1PHIHn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L1PHIHn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L1PHIHn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L1PHIHn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L1PHIHn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L1PHIHn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L1PHIHn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L1PHIHn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L1PHIHn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L1PHIHn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L1PHIHn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L1PHIHn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L1PHIHn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L1PHIHn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L1PHIHn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L1PHIHn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L1PHIHn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L1PHIHn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L1PHIHn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L1PHIHn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L1PHIHn2_enb,
      allstub_dataarray_data_V_address0  => AS_L1PHIHn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L1PHIHn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L1PHIH_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L1PHIH_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L1PHIH_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L1PHIH_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L1PHIH_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L1PHIH_din
  );

  LATCH_MP_L2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L2PHIA_bx,
      start => MP_L2PHIA_start
  );

  MP_L2PHIA : entity work.MP_L2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L2PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L2PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L3L4AB_L2PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L3L4AB_L2PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L3L4AB_L2PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L3L4AB_L2PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L3L4AB_L2PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L2PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L2PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L5L6ABCD_L2PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L5L6ABCD_L2PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L5L6ABCD_L2PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L2PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L2PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_D1D2ABCD_L2PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_D1D2ABCD_L2PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_D1D2ABCD_L2PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L2PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L2PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L2PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L2PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L2PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L2PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L2PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L2PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L2PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L2PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L2PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L2PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L2PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L2PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L2PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L2PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L2PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L2PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L2PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L2PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L2PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L2PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L2PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L2PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L2PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L2PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L2PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L2PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L2PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L2PHIA_din
  );

  LATCH_MP_L2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L2PHIB_bx,
      start => MP_L2PHIB_start
  );

  MP_L2PHIB : entity work.MP_L2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L2PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L2PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L3L4AB_L2PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L3L4AB_L2PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L3L4AB_L2PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L3L4AB_L2PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L3L4AB_L2PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4CD_L2PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4CD_L2PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4CD_L2PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4CD_L2PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4CD_L2PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L2PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L2PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L2PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L2PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L2PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L2PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L2PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L2PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L2PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L2PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L2PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L2PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L2PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L2PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L2PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L2PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L2PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L2PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L2PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L2PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L2PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L2PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L2PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L2PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L2PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L2PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L2PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L2PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L2PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L2PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L2PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L2PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L2PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L2PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L2PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L2PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L2PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L2PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L2PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L2PHIB_din
  );

  LATCH_MP_L2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L2PHIC_bx,
      start => MP_L2PHIC_start
  );

  MP_L2PHIC : entity work.MP_L2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L2PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L2PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L3L4AB_L2PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L3L4AB_L2PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L3L4AB_L2PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L3L4AB_L2PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L3L4AB_L2PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L3L4AB_L2PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L3L4CD_L2PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L3L4CD_L2PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L3L4CD_L2PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L3L4CD_L2PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L3L4CD_L2PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L2PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L2PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L2PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L2PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L2PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L2PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L2PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_D1D2ABCD_L2PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_D1D2ABCD_L2PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_D1D2ABCD_L2PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L2PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L2PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L2PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L2PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L2PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L2PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L2PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L2PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L2PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L2PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L2PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L2PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L2PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L2PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L2PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L2PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L2PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L2PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L2PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L2PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L2PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L2PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L2PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L2PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L2PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L2PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L2PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L2PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L2PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L2PHIC_din
  );

  LATCH_MP_L2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L2PHID_bx,
      start => MP_L2PHID_start
  );

  MP_L2PHID : entity work.MP_L2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L2PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L2PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L3L4CD_L2PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L3L4CD_L2PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L3L4CD_L2PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L3L4CD_L2PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L3L4CD_L2PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L3L4CD_L2PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L2PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L2PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L2PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L5L6ABCD_L2PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L5L6ABCD_L2PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L5L6ABCD_L2PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_L2PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_D1D2ABCD_L2PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_D1D2ABCD_L2PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_D1D2ABCD_L2PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_D1D2ABCD_L2PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_D1D2ABCD_L2PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L2PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L2PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L2PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L2PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L2PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L2PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L2PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L2PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L2PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L2PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L2PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L2PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L2PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L2PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L2PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L2PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L2PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L2PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L2PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L2PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L2PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L2PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L2PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L2PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L2PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L2PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L2PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L2PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L2PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L2PHID_din
  );

  LATCH_MP_L3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L3PHIA_bx,
      start => MP_L3PHIA_start
  );

  MP_L3PHIA : entity work.MP_L3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L3PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L3PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L3PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L3PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L3PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L3PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L3PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L3PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L3PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L3PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L3PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L3PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L3PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L3PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L3PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L3PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L3PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L3PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L3PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L3PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L3PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L3PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L3PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L3PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L3PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L3PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L3PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L3PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L3PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L3PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L3PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L3PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L3PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L3PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L3PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L3PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L3PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L3PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L3PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L3PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L3PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L3PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L3PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L3PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L3PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L3PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L3PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L3PHIA_din
  );

  LATCH_MP_L3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L3PHIB_bx,
      start => MP_L3PHIB_start
  );

  MP_L3PHIB : entity work.MP_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L3PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L3PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L3PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L3PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L3PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L3PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L3PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L3PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L3PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L3PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L3PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L3PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L3PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L3PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L3PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L3PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L3PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L3PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L3PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_L3PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_L3PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_L3PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_L3PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_L3PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_L3PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_L3PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_L3PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_L3PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_L3PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_L3PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L3PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L3PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L5L6ABCD_L3PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L5L6ABCD_L3PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L5L6ABCD_L3PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L3PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L3PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L3PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L3PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L3PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L3PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L3PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L3PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L3PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L3PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L3PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L3PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L3PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L3PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L3PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L3PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L3PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L3PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L3PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L3PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L3PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L3PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L3PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L3PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L3PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L3PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L3PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L3PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L3PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L3PHIB_din
  );

  LATCH_MP_L3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L3PHIC_bx,
      start => MP_L3PHIC_start
  );

  MP_L3PHIC : entity work.MP_L3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L3PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L3PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_L3PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_L3PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_L3PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_L3PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_L3PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_L3PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_L3PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_L3PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_L3PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_L3PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_L3PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_L3PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_L3PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_L3PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_L3PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_L3PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_L3PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_L3PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_L3PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_L3PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_L3PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_L3PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_L3PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L3PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_L3PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_L3PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_L3PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_L3PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_L3PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L3PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L3PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L5L6ABCD_L3PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L5L6ABCD_L3PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L5L6ABCD_L3PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L3PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L3PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L3PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L3PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L3PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L3PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L3PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L3PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L3PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L3PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L3PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L3PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L3PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L3PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L3PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L3PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L3PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L3PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L3PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L3PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L3PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L3PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L3PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L3PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L3PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L3PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L3PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L3PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L3PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L3PHIC_din
  );

  LATCH_MP_L3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L3PHID_bx,
      start => MP_L3PHID_start
  );

  MP_L3PHID : entity work.MP_L3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L3PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L3PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2HI_L3PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2HI_L3PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2HI_L3PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2HI_L3PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2HI_L3PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2HI_L3PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L3PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2JKL_L3PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2JKL_L3PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2JKL_L3PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2JKL_L3PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2JKL_L3PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L3PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L3PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L3PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L5L6ABCD_L3PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L5L6ABCD_L3PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L5L6ABCD_L3PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L3PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L3PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L3PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L3PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L3PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L3PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L3PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L3PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L3PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L3PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L3PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L3PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L3PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L3PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L3PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L3PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L3PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L3PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L3PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L3PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L3PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L3PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L3PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L3PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L3PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L3PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L3PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L3PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L3PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L3PHID_din
  );

  LATCH_MP_L4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L4PHIA_bx,
      start => MP_L4PHIA_start
  );

  MP_L4PHIA : entity work.MP_L4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L4PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L4PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L4PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L4PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L4PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L4PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L4PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L4PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L4PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L4PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L4PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L4PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L4PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L4PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L4PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L4PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L4PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L4PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L4PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L4PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_L4PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_L4PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_L4PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L4PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L4PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_L5L6ABCD_L4PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L5L6ABCD_L4PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L5L6ABCD_L4PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L4PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L4PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L4PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L4PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L4PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L4PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L4PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L4PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L4PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L4PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L4PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L4PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L4PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L4PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L4PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L4PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L4PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L4PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L4PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L4PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L4PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L4PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L4PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L4PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L4PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L4PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L4PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L4PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L4PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L4PHIA_din
  );

  LATCH_MP_L4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L4PHIB_bx,
      start => MP_L4PHIB_start
  );

  MP_L4PHIB : entity work.MP_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L4PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L4PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L4PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L4PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L4PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L4PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L4PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L4PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L4PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L4PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L4PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L4PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L4PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L4PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L4PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L4PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L4PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L4PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_L4PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_L4PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_L4PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_L4PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_L4PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_L4PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_L4PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_L4PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_L4PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_L4PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L4PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L4PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_L4PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_L4PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_L4PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L4PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L4PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_L5L6ABCD_L4PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L5L6ABCD_L4PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L5L6ABCD_L4PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L4PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L4PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L4PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L4PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L4PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L4PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L4PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L4PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L4PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L4PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L4PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L4PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L4PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L4PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L4PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L4PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L4PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L4PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L4PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L4PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L4PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L4PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L4PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L4PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L4PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L4PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L4PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L4PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L4PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L4PHIB_din
  );

  LATCH_MP_L4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L4PHIC_bx,
      start => MP_L4PHIC_start
  );

  MP_L4PHIC : entity work.MP_L4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L4PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L4PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_L4PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_L4PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_L4PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_L4PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_L4PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_L4PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_L4PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_L4PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_L4PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_L4PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_L4PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_L4PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_L4PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_L4PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_L4PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_L4PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_L4PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_L4PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_L4PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_L4PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_L4PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_L4PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L4PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_L4PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_L4PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_L4PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_L4PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_L4PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L4PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L4PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_L4PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_L4PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_L4PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L4PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L4PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_L5L6ABCD_L4PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L5L6ABCD_L4PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L5L6ABCD_L4PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L4PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L4PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L4PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L4PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L4PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L4PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L4PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L4PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L4PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L4PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L4PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L4PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L4PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L4PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L4PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L4PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L4PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L4PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L4PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L4PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L4PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L4PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L4PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L4PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L4PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L4PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L4PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L4PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L4PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L4PHIC_din
  );

  LATCH_MP_L4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L4PHID_bx,
      start => MP_L4PHID_start
  );

  MP_L4PHID : entity work.MP_L4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L4PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L4PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_L4PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_L4PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_L4PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_L4PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_L4PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_L4PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_L4PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_L4PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_L4PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_L4PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_L4PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_L4PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L4PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_L4PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_L4PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_L4PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_L4PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_L4PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L4PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L4PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L4PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_L4PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_L4PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_L4PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L5L6ABCD_L4PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L5L6ABCD_L4PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L5L6ABCD_L4PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_L5L6ABCD_L4PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L5L6ABCD_L4PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L5L6ABCD_L4PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L4PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L4PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L4PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L4PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L4PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L4PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L4PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L4PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L4PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L4PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L4PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L4PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L4PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L4PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L4PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L4PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L4PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L4PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L4PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L4PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L4PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L4PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L4PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L4PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L4PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L4PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L4PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L4PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L4PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L4PHID_din
  );

  LATCH_MP_L5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L5PHIA_bx,
      start => MP_L5PHIA_start
  );

  MP_L5PHIA : entity work.MP_L5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L5PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L5PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L5PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L5PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L5PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L5PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L5PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L5PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L5PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L5PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L5PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L5PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L5PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L5PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L5PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L5PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L5PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L5PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L5PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L5PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_L5PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_L5PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_L5PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4AB_L5PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4AB_L5PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4AB_L5PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4AB_L5PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4AB_L5PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L5PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L5PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L5PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L5PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L5PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L5PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L5PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L5PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L5PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L5PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L5PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L5PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L5PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L5PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L5PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L5PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L5PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L5PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L5PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L5PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L5PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L5PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L5PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L5PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L5PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L5PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L5PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L5PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L5PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L5PHIA_din
  );

  LATCH_MP_L5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L5PHIB_bx,
      start => MP_L5PHIB_start
  );

  MP_L5PHIB : entity work.MP_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L5PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L5PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L5PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L5PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L5PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L5PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L5PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L5PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L5PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L5PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L5PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L5PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L5PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L5PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L5PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L5PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L5PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L5PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_L5PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_L5PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_L5PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_L5PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_L5PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_L5PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_L5PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_L5PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_L5PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_L5PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L5PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L5PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_L5PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_L5PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_L5PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_L5PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_L5PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_L5PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_L5PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_L5PHIB_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_L5PHIB_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHIB_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_L5PHIB_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_L5PHIB_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_L5PHIB_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_L5PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L5PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L5PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L5PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L5PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L5PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L5PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L5PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L5PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L5PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L5PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L5PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L5PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L5PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L5PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L5PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L5PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L5PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L5PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L5PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L5PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L5PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L5PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L5PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L5PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L5PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L5PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L5PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L5PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L5PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L5PHIB_din
  );

  LATCH_MP_L5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L5PHIC_bx,
      start => MP_L5PHIC_start
  );

  MP_L5PHIC : entity work.MP_L5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L5PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L5PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_L5PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_L5PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_L5PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_L5PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_L5PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_L5PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_L5PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_L5PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_L5PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_L5PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_L5PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_L5PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_L5PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_L5PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_L5PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_L5PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_L5PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_L5PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_L5PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_L5PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_L5PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_L5PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L5PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_L5PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_L5PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_L5PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_L5PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_L5PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L5PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L5PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_L5PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_L5PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_L5PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_L5PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_L5PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_L5PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_L5PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_L5PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_L5PHIC_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_L5PHIC_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHIC_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_L5PHIC_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_L5PHIC_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_L5PHIC_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_L5PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L5PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L5PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L5PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L5PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L5PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L5PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L5PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L5PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L5PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L5PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L5PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L5PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L5PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L5PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L5PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L5PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L5PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L5PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L5PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L5PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L5PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L5PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L5PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L5PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L5PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L5PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L5PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L5PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L5PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L5PHIC_din
  );

  LATCH_MP_L5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L5PHID_bx,
      start => MP_L5PHID_start
  );

  MP_L5PHID : entity work.MP_L5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L5PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L5PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_L5PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_L5PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_L5PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_L5PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_L5PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_L5PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_L5PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_L5PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_L5PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_L5PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_L5PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_L5PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L5PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_L5PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_L5PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_L5PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_L5PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_L5PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_L5PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_L5PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_L5PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_L5PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_L5PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_L5PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4CD_L5PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4CD_L5PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4CD_L5PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4CD_L5PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4CD_L5PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4CD_L5PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L5PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L5PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L5PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L5PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L5PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L5PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L5PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L5PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L5PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L5PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L5PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L5PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L5PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L5PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L5PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L5PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L5PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L5PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L5PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L5PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L5PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L5PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L5PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L5PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L5PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L5PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L5PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L5PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L5PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L5PHID_din
  );

  LATCH_MP_L6PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L6PHIA_bx,
      start => MP_L6PHIA_start
  );

  MP_L6PHIA : entity work.MP_L6PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L6PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L6PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L6PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L6PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L6PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L6PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L6PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L6PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L6PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L6PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L6PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L6PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L6PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L6PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L6PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L6PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L6PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L6PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L3L4AB_L6PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L3L4AB_L6PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L3L4AB_L6PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L3L4AB_L6PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L3L4AB_L6PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L6PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L6PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L6PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L6PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L6PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L6PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L6PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L6PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L6PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L6PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L6PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L6PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L6PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L6PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L6PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L6PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L6PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L6PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L6PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L6PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L6PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L6PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_L6PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L6PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L6PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L6PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L6PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L6PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L6PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L6PHIA_din
  );

  LATCH_MP_L6PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L6PHIB_bx,
      start => MP_L6PHIB_start
  );

  MP_L6PHIB : entity work.MP_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L6PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L6PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_L6PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_L6PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_L6PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_L6PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_L6PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_L6PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_L6PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_L6PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_L6PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_L6PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_L6PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_L6PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_L6PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_L6PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_L6PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_L6PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_L6PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_L6PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_L6PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_L6PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_L6PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_L6PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_L6PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_L6PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_L6PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_L6PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L3L4AB_L6PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L3L4AB_L6PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L3L4AB_L6PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L3L4AB_L6PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L3L4AB_L6PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4CD_L6PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4CD_L6PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4CD_L6PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4CD_L6PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4CD_L6PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L6PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L6PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L6PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L6PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L6PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L6PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L6PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L6PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L6PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L6PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L6PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L6PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L6PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L6PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L6PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L6PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L6PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L6PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L6PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L6PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L6PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L6PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_L6PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L6PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L6PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L6PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L6PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L6PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L6PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L6PHIB_din
  );

  LATCH_MP_L6PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L6PHIC_bx,
      start => MP_L6PHIC_start
  );

  MP_L6PHIC : entity work.MP_L6PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L6PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L6PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_L6PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_L6PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_L6PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_L6PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_L6PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_L6PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_L6PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_L6PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_L6PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_L6PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_L6PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_L6PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_L6PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_L6PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_L6PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_L6PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_L6PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_L6PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_L6PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_L6PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_L6PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_L6PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L6PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_L6PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_L6PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_L6PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_L6PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_L6PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L3L4AB_L6PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L3L4AB_L6PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L3L4AB_L6PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L3L4AB_L6PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L3L4AB_L6PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L3L4AB_L6PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4CD_L6PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4CD_L6PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4CD_L6PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4CD_L6PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4CD_L6PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L6PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L6PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L6PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L6PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L6PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L6PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L6PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L6PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L6PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L6PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L6PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L6PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L6PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L6PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L6PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L6PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L6PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L6PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L6PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L6PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L6PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L6PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_L6PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L6PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L6PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L6PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L6PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L6PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L6PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L6PHIC_din
  );

  LATCH_MP_L6PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_L6PHID_bx,
      start => MP_L6PHID_start
  );

  MP_L6PHID : entity work.MP_L6PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_L6PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_L6PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_L6PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_L6PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_L6PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_L6PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_L6PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_L6PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_L6PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_L6PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_L6PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_L6PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_L6PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_L6PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_L6PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_L6PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_L6PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_L6PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_L6PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_L6PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L3L4CD_L6PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L3L4CD_L6PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L3L4CD_L6PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L3L4CD_L6PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L3L4CD_L6PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L3L4CD_L6PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_L6PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_L6PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_L6PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_L6PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_L6PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_L6PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_L6PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_L6PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_L6PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_L6PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_L6PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_L6PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_L6PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_L6PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_L6PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_L6PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_L6PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_L6PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_L6PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_L6PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_L6PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_L6PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_L6PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_L6PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_L6PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_L6PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_L6PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_L6PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_L6PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_L6PHID_din
  );

  LATCH_MP_D1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D1PHIA_bx,
      start => MP_D1PHIA_start
  );

  MP_D1PHIA : entity work.MP_D1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D1PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D1PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D1PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D1PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D1PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D1PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D1PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D1PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D1PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D1PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D1PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D1PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D1PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D1PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D1PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D1PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D1PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D1PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D1PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D1PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D1PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D1PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D1PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4AB_D1PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4AB_D1PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4AB_D1PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4AB_D1PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4AB_D1PHIA_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D1PHIA_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIA_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D1PHIA_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_D1PHIA_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_D1PHIA_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_D1PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D1PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D1PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D1PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D1PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D1PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D1PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D1PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D1PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D1PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D1PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D1PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D1PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D1PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D1PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D1PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D1PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D1PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D1PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D1PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D1PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D1PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D1PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_D1PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D1PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D1PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D1PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D1PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D1PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D1PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D1PHIA_din
  );

  LATCH_MP_D1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D1PHIB_bx,
      start => MP_D1PHIB_start
  );

  MP_D1PHIB : entity work.MP_D1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D1PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D1PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D1PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D1PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D1PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D1PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D1PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D1PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D1PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D1PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D1PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D1PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D1PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D1PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D1PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D1PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D1PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D1PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_D1PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_D1PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_D1PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_D1PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_D1PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_D1PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_D1PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_D1PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_D1PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_D1PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D1PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D1PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D1PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D1PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D1PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_D1PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_D1PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_D1PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_D1PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_D1PHIB_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_D1PHIB_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHIB_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_D1PHIB_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_D1PHIB_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_D1PHIB_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_D1PHIB_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D1PHIB_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIB_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D1PHIB_V_dout,
      projin_8_mask_0_V                   => MPROJ_D3D4ABCD_D1PHIB_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_D3D4ABCD_D1PHIB_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_D3D4ABCD_D1PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D1PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D1PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D1PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D1PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D1PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D1PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D1PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D1PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D1PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D1PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D1PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D1PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D1PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D1PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D1PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D1PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D1PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D1PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D1PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D1PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D1PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D1PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_D1PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D1PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D1PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D1PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D1PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D1PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D1PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D1PHIB_din
  );

  LATCH_MP_D1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D1PHIC_bx,
      start => MP_D1PHIC_start
  );

  MP_D1PHIC : entity work.MP_D1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D1PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D1PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_D1PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_D1PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_D1PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_D1PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_D1PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_D1PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_D1PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_D1PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_D1PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_D1PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_D1PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_D1PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_D1PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_D1PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_D1PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_D1PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_D1PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_D1PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_D1PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_D1PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_D1PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_D1PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D1PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_D1PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_D1PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_D1PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_D1PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_D1PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D1PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D1PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D1PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D1PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D1PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_D1PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_D1PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_D1PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_D1PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_D1PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_D1PHIC_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_D1PHIC_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHIC_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_D1PHIC_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_D1PHIC_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_D1PHIC_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_D1PHIC_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D1PHIC_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHIC_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D1PHIC_V_dout,
      projin_8_mask_0_V                   => MPROJ_D3D4ABCD_D1PHIC_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_D3D4ABCD_D1PHIC_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_D3D4ABCD_D1PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D1PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D1PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D1PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D1PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D1PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D1PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D1PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D1PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D1PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D1PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D1PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D1PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D1PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D1PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D1PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D1PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D1PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D1PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D1PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D1PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D1PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D1PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_D1PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D1PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D1PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D1PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D1PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D1PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D1PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D1PHIC_din
  );

  LATCH_MP_D1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D1PHID_bx,
      start => MP_D1PHID_start
  );

  MP_D1PHID : entity work.MP_D1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D1PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D1PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_D1PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_D1PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_D1PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_D1PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_D1PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_D1PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_D1PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_D1PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_D1PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_D1PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_D1PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_D1PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D1PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_D1PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_D1PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_D1PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_D1PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_D1PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D1PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D1PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D1PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D1PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D1PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D1PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4CD_D1PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4CD_D1PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4CD_D1PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4CD_D1PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4CD_D1PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4CD_D1PHID_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D1PHID_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D1PHID_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D1PHID_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_D1PHID_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_D1PHID_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_D1PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D1PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D1PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D1PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D1PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D1PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D1PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D1PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D1PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D1PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D1PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D1PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D1PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D1PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D1PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D1PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D1PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D1PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D1PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D1PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D1PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D1PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D1PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_D1PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D1PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D1PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D1PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D1PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D1PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D1PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D1PHID_din
  );

  LATCH_MP_D2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D2PHIA_bx,
      start => MP_D2PHIA_start
  );

  MP_D2PHIA : entity work.MP_D2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D2PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D2PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D2PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D2PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D2PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D2PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D2PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D2PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D2PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D2PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D2PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D2PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D2PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D2PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D2PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D2PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D2PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D2PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D2PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D2PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D2PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D2PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D2PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4AB_D2PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4AB_D2PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4AB_D2PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4AB_D2PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4AB_D2PHIA_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D2PHIA_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIA_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D2PHIA_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_D2PHIA_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_D2PHIA_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_D2PHIA_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D2PHIA_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIA_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D2PHIA_V_dout,
      projin_6_mask_0_V                   => MPROJ_L1D1ABCD_D2PHIA_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L1D1ABCD_D2PHIA_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L1D1ABCD_D2PHIA_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D2PHIA_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIA_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D2PHIA_V_dout,
      projin_7_mask_0_V                   => MPROJ_L2D1ABCD_D2PHIA_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L2D1ABCD_D2PHIA_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L2D1ABCD_D2PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D2PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D2PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D2PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D2PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D2PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D2PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D2PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D2PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D2PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D2PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D2PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D2PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D2PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D2PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D2PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D2PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D2PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D2PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D2PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D2PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D2PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D2PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_D2PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D2PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D2PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D2PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D2PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D2PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D2PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D2PHIA_din
  );

  LATCH_MP_D2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D2PHIB_bx,
      start => MP_D2PHIB_start
  );

  MP_D2PHIB : entity work.MP_D2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D2PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D2PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D2PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D2PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D2PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D2PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D2PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D2PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D2PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D2PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D2PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D2PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D2PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D2PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D2PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D2PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D2PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D2PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_D2PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_D2PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_D2PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_D2PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_D2PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_D2PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_D2PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_D2PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_D2PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_D2PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D2PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D2PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D2PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D2PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D2PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_D2PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_D2PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_D2PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_D2PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_D2PHIB_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_D2PHIB_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHIB_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_D2PHIB_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_D2PHIB_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_D2PHIB_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_D2PHIB_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D2PHIB_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIB_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D2PHIB_V_dout,
      projin_8_mask_0_V                   => MPROJ_D3D4ABCD_D2PHIB_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_D3D4ABCD_D2PHIB_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_D3D4ABCD_D2PHIB_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D2PHIB_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIB_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D2PHIB_V_dout,
      projin_9_mask_0_V                   => MPROJ_L1D1ABCD_D2PHIB_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L1D1ABCD_D2PHIB_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L1D1ABCD_D2PHIB_AV_dout_nent(7),
      projin_10_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D2PHIB_enb,
      projin_10_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHIB_V_readaddr,
      projin_10_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D2PHIB_V_dout,
      projin_10_mask_0_V                   => MPROJ_L1D1EFGH_D2PHIB_AV_dout_mask(0),
      projin_10_mask_1_V                   => MPROJ_L1D1EFGH_D2PHIB_AV_dout_mask(1),
      projin_10_nentries_0_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(0),
      projin_10_nentries_1_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(1),
      projin_10_nentries_2_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(2),
      projin_10_nentries_3_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(3),
      projin_10_nentries_4_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(4),
      projin_10_nentries_5_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(5),
      projin_10_nentries_6_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(6),
      projin_10_nentries_7_V               => MPROJ_L1D1EFGH_D2PHIB_AV_dout_nent(7),
      projin_11_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D2PHIB_enb,
      projin_11_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIB_V_readaddr,
      projin_11_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D2PHIB_V_dout,
      projin_11_mask_0_V                   => MPROJ_L2D1ABCD_D2PHIB_AV_dout_mask(0),
      projin_11_mask_1_V                   => MPROJ_L2D1ABCD_D2PHIB_AV_dout_mask(1),
      projin_11_nentries_0_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(0),
      projin_11_nentries_1_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(1),
      projin_11_nentries_2_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(2),
      projin_11_nentries_3_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(3),
      projin_11_nentries_4_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(4),
      projin_11_nentries_5_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(5),
      projin_11_nentries_6_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(6),
      projin_11_nentries_7_V               => MPROJ_L2D1ABCD_D2PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D2PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D2PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D2PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D2PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D2PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D2PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D2PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D2PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D2PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D2PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D2PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D2PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D2PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D2PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D2PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D2PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D2PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D2PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D2PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D2PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D2PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D2PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_D2PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D2PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D2PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D2PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D2PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D2PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D2PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D2PHIB_din
  );

  LATCH_MP_D2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D2PHIC_bx,
      start => MP_D2PHIC_start
  );

  MP_D2PHIC : entity work.MP_D2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D2PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D2PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_D2PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_D2PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_D2PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_D2PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_D2PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_D2PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_D2PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_D2PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_D2PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_D2PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_D2PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_D2PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_D2PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_D2PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_D2PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_D2PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_D2PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_D2PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_D2PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_D2PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_D2PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_D2PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D2PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_D2PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_D2PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_D2PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_D2PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_D2PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D2PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D2PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D2PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D2PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D2PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L3L4AB_D2PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L3L4AB_D2PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L3L4AB_D2PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_L3L4AB_D2PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L3L4AB_D2PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L3L4AB_D2PHIC_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L3L4CD_D2PHIC_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHIC_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L3L4CD_D2PHIC_V_dout,
      projin_7_mask_0_V                   => MPROJ_L3L4CD_D2PHIC_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L3L4CD_D2PHIC_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L3L4CD_D2PHIC_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D2PHIC_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHIC_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D2PHIC_V_dout,
      projin_8_mask_0_V                   => MPROJ_D3D4ABCD_D2PHIC_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_D3D4ABCD_D2PHIC_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_D3D4ABCD_D2PHIC_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D2PHIC_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D2PHIC_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D2PHIC_V_dout,
      projin_9_mask_0_V                   => MPROJ_L1D1ABCD_D2PHIC_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L1D1ABCD_D2PHIC_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L1D1ABCD_D2PHIC_AV_dout_nent(7),
      projin_10_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D2PHIC_enb,
      projin_10_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHIC_V_readaddr,
      projin_10_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D2PHIC_V_dout,
      projin_10_mask_0_V                   => MPROJ_L1D1EFGH_D2PHIC_AV_dout_mask(0),
      projin_10_mask_1_V                   => MPROJ_L1D1EFGH_D2PHIC_AV_dout_mask(1),
      projin_10_nentries_0_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(0),
      projin_10_nentries_1_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(1),
      projin_10_nentries_2_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(2),
      projin_10_nentries_3_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(3),
      projin_10_nentries_4_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(4),
      projin_10_nentries_5_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(5),
      projin_10_nentries_6_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(6),
      projin_10_nentries_7_V               => MPROJ_L1D1EFGH_D2PHIC_AV_dout_nent(7),
      projin_11_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D2PHIC_enb,
      projin_11_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHIC_V_readaddr,
      projin_11_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D2PHIC_V_dout,
      projin_11_mask_0_V                   => MPROJ_L2D1ABCD_D2PHIC_AV_dout_mask(0),
      projin_11_mask_1_V                   => MPROJ_L2D1ABCD_D2PHIC_AV_dout_mask(1),
      projin_11_nentries_0_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(0),
      projin_11_nentries_1_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(1),
      projin_11_nentries_2_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(2),
      projin_11_nentries_3_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(3),
      projin_11_nentries_4_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(4),
      projin_11_nentries_5_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(5),
      projin_11_nentries_6_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(6),
      projin_11_nentries_7_V               => MPROJ_L2D1ABCD_D2PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D2PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D2PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D2PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D2PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D2PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D2PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D2PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D2PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D2PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D2PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D2PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D2PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D2PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D2PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D2PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D2PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D2PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D2PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D2PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D2PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D2PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D2PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_D2PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D2PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D2PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D2PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D2PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D2PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D2PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D2PHIC_din
  );

  LATCH_MP_D2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D2PHID_bx,
      start => MP_D2PHID_start
  );

  MP_D2PHID : entity work.MP_D2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D2PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D2PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_D2PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_D2PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_D2PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_D2PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_D2PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_D2PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_D2PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_D2PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_D2PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_D2PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_D2PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_D2PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D2PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_D2PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_D2PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_D2PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_D2PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_D2PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D2PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D2PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D2PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D2PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D2PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D2PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L3L4CD_D2PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L3L4CD_D2PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L3L4CD_D2PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_L3L4CD_D2PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L3L4CD_D2PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L3L4CD_D2PHID_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D2PHID_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D2PHID_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D2PHID_V_dout,
      projin_5_mask_0_V                   => MPROJ_D3D4ABCD_D2PHID_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_D3D4ABCD_D2PHID_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_D3D4ABCD_D2PHID_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D2PHID_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D2PHID_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D2PHID_V_dout,
      projin_6_mask_0_V                   => MPROJ_L1D1EFGH_D2PHID_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L1D1EFGH_D2PHID_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L1D1EFGH_D2PHID_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D2PHID_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D2PHID_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D2PHID_V_dout,
      projin_7_mask_0_V                   => MPROJ_L2D1ABCD_D2PHID_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L2D1ABCD_D2PHID_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L2D1ABCD_D2PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D2PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D2PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D2PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D2PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D2PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D2PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D2PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D2PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D2PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D2PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D2PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D2PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D2PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D2PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D2PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D2PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D2PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D2PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D2PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D2PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D2PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D2PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_D2PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D2PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D2PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D2PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D2PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D2PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D2PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D2PHID_din
  );

  LATCH_MP_D3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D3PHIA_bx,
      start => MP_D3PHIA_start
  );

  MP_D3PHIA : entity work.MP_D3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D3PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D3PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D3PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D3PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D3PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D3PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D3PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D3PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D3PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D3PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D3PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D3PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D3PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D3PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D3PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D3PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D3PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D3PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D3PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D3PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D3PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D3PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D3PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D3PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D3PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_D3PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_D3PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_D3PHIA_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D3PHIA_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIA_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D3PHIA_V_dout,
      projin_5_mask_0_V                   => MPROJ_L1D1ABCD_D3PHIA_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L1D1ABCD_D3PHIA_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L1D1ABCD_D3PHIA_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D3PHIA_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIA_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D3PHIA_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_D3PHIA_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_D3PHIA_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_D3PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D3PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D3PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D3PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D3PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D3PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D3PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D3PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D3PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D3PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D3PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D3PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D3PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D3PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D3PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D3PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D3PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D3PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D3PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D3PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D3PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D3PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D3PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_D3PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D3PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D3PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D3PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D3PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D3PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D3PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D3PHIA_din
  );

  LATCH_MP_D3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D3PHIB_bx,
      start => MP_D3PHIB_start
  );

  MP_D3PHIB : entity work.MP_D3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D3PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D3PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D3PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D3PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D3PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D3PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D3PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D3PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D3PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D3PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D3PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D3PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D3PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D3PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D3PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D3PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D3PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D3PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_D3PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_D3PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_D3PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_D3PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_D3PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_D3PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_D3PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_D3PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_D3PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_D3PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D3PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D3PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D3PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D3PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D3PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D3PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D3PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_D1D2ABCD_D3PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_D1D2ABCD_D3PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_D1D2ABCD_D3PHIB_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D3PHIB_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIB_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D3PHIB_V_dout,
      projin_7_mask_0_V                   => MPROJ_L1D1ABCD_D3PHIB_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L1D1ABCD_D3PHIB_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L1D1ABCD_D3PHIB_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D3PHIB_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHIB_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D3PHIB_V_dout,
      projin_8_mask_0_V                   => MPROJ_L1D1EFGH_D3PHIB_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_L1D1EFGH_D3PHIB_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_L1D1EFGH_D3PHIB_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D3PHIB_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIB_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D3PHIB_V_dout,
      projin_9_mask_0_V                   => MPROJ_L2D1ABCD_D3PHIB_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L2D1ABCD_D3PHIB_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L2D1ABCD_D3PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D3PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D3PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D3PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D3PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D3PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D3PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D3PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D3PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D3PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D3PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D3PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D3PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D3PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D3PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D3PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D3PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D3PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D3PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D3PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D3PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D3PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D3PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_D3PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D3PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D3PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D3PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D3PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D3PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D3PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D3PHIB_din
  );

  LATCH_MP_D3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D3PHIC_bx,
      start => MP_D3PHIC_start
  );

  MP_D3PHIC : entity work.MP_D3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D3PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D3PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_D3PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_D3PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_D3PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_D3PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_D3PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_D3PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_D3PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_D3PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_D3PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_D3PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_D3PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_D3PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_D3PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_D3PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_D3PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_D3PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_D3PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_D3PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_D3PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_D3PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_D3PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_D3PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D3PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_D3PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_D3PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_D3PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_D3PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_D3PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D3PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D3PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D3PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D3PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D3PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D3PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D3PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_D1D2ABCD_D3PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_D1D2ABCD_D3PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_D1D2ABCD_D3PHIC_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D3PHIC_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D3PHIC_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D3PHIC_V_dout,
      projin_7_mask_0_V                   => MPROJ_L1D1ABCD_D3PHIC_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L1D1ABCD_D3PHIC_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L1D1ABCD_D3PHIC_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D3PHIC_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHIC_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D3PHIC_V_dout,
      projin_8_mask_0_V                   => MPROJ_L1D1EFGH_D3PHIC_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_L1D1EFGH_D3PHIC_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_L1D1EFGH_D3PHIC_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D3PHIC_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHIC_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D3PHIC_V_dout,
      projin_9_mask_0_V                   => MPROJ_L2D1ABCD_D3PHIC_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L2D1ABCD_D3PHIC_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L2D1ABCD_D3PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D3PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D3PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D3PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D3PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D3PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D3PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D3PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D3PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D3PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D3PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D3PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D3PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D3PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D3PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D3PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D3PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D3PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D3PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D3PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D3PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D3PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D3PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_D3PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D3PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D3PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D3PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D3PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D3PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D3PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D3PHIC_din
  );

  LATCH_MP_D3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D3PHID_bx,
      start => MP_D3PHID_start
  );

  MP_D3PHID : entity work.MP_D3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D3PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D3PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_D3PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_D3PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_D3PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_D3PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_D3PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_D3PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_D3PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_D3PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_D3PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_D3PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_D3PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_D3PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D3PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_D3PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_D3PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_D3PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_D3PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_D3PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D3PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D3PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D3PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D3PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D3PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D3PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D3PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D3PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D3PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_D3PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_D3PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_D3PHID_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D3PHID_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D3PHID_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D3PHID_V_dout,
      projin_5_mask_0_V                   => MPROJ_L1D1EFGH_D3PHID_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L1D1EFGH_D3PHID_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L1D1EFGH_D3PHID_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D3PHID_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D3PHID_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D3PHID_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_D3PHID_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_D3PHID_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_D3PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D3PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D3PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D3PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D3PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D3PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D3PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D3PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D3PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D3PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D3PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D3PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D3PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D3PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D3PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D3PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D3PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D3PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D3PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D3PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D3PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D3PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D3PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_D3PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D3PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D3PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D3PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D3PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D3PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D3PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D3PHID_din
  );

  LATCH_MP_D4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D4PHIA_bx,
      start => MP_D4PHIA_start
  );

  MP_D4PHIA : entity work.MP_D4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D4PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D4PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D4PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D4PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D4PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D4PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D4PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D4PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D4PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D4PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D4PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D4PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D4PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D4PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D4PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D4PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D4PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D4PHIA_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D4PHIA_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIA_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D4PHIA_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D4PHIA_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D4PHIA_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D4PHIA_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D4PHIA_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIA_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D4PHIA_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_D4PHIA_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_D4PHIA_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_D4PHIA_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D4PHIA_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIA_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D4PHIA_V_dout,
      projin_5_mask_0_V                   => MPROJ_L1D1ABCD_D4PHIA_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L1D1ABCD_D4PHIA_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L1D1ABCD_D4PHIA_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D4PHIA_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIA_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D4PHIA_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_D4PHIA_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_D4PHIA_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_D4PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D4PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D4PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D4PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D4PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D4PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D4PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D4PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D4PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D4PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D4PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D4PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D4PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D4PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D4PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D4PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D4PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D4PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D4PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D4PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D4PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D4PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D4PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_D4PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D4PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D4PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D4PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D4PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D4PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D4PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D4PHIA_din
  );

  LATCH_MP_D4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D4PHIB_bx,
      start => MP_D4PHIB_start
  );

  MP_D4PHIB : entity work.MP_D4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D4PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D4PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2ABC_D4PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2ABC_D4PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2ABC_D4PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2ABC_D4PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2ABC_D4PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2ABC_D4PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2DE_D4PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2DE_D4PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2DE_D4PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2DE_D4PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2DE_D4PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2F_D4PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2F_D4PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2F_D4PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2F_D4PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2F_D4PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2G_D4PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2G_D4PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2G_D4PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2G_D4PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2G_D4PHIB_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2HI_D4PHIB_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHIB_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2HI_D4PHIB_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2HI_D4PHIB_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2HI_D4PHIB_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2HI_D4PHIB_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D4PHIB_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIB_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D4PHIB_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D4PHIB_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D4PHIB_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D4PHIB_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D4PHIB_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIB_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D4PHIB_V_dout,
      projin_6_mask_0_V                   => MPROJ_D1D2ABCD_D4PHIB_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_D1D2ABCD_D4PHIB_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_D1D2ABCD_D4PHIB_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D4PHIB_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIB_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D4PHIB_V_dout,
      projin_7_mask_0_V                   => MPROJ_L1D1ABCD_D4PHIB_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L1D1ABCD_D4PHIB_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L1D1ABCD_D4PHIB_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D4PHIB_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHIB_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D4PHIB_V_dout,
      projin_8_mask_0_V                   => MPROJ_L1D1EFGH_D4PHIB_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_L1D1EFGH_D4PHIB_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_L1D1EFGH_D4PHIB_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D4PHIB_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIB_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D4PHIB_V_dout,
      projin_9_mask_0_V                   => MPROJ_L2D1ABCD_D4PHIB_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L2D1ABCD_D4PHIB_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L2D1ABCD_D4PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D4PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D4PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D4PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D4PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D4PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D4PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D4PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D4PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D4PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D4PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D4PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D4PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D4PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D4PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D4PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D4PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D4PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D4PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D4PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D4PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D4PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D4PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_D4PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D4PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D4PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D4PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D4PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D4PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D4PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D4PHIB_din
  );

  LATCH_MP_D4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D4PHIC_bx,
      start => MP_D4PHIC_start
  );

  MP_D4PHIC : entity work.MP_D4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D4PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D4PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2DE_D4PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2DE_D4PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2DE_D4PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2DE_D4PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2DE_D4PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2DE_D4PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2F_D4PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2F_D4PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2F_D4PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2F_D4PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2F_D4PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2F_D4PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2G_D4PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2G_D4PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2G_D4PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2G_D4PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2G_D4PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1L2HI_D4PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1L2HI_D4PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1L2HI_D4PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1L2HI_D4PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1L2HI_D4PHIC_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D4PHIC_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_L1L2JKL_D4PHIC_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_L1L2JKL_D4PHIC_V_dout,
      projin_4_mask_0_V                   => MPROJ_L1L2JKL_D4PHIC_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_L1L2JKL_D4PHIC_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_L1L2JKL_D4PHIC_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D4PHIC_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHIC_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D4PHIC_V_dout,
      projin_5_mask_0_V                   => MPROJ_L2L3ABCD_D4PHIC_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L2L3ABCD_D4PHIC_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L2L3ABCD_D4PHIC_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D4PHIC_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHIC_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D4PHIC_V_dout,
      projin_6_mask_0_V                   => MPROJ_D1D2ABCD_D4PHIC_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_D1D2ABCD_D4PHIC_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_D1D2ABCD_D4PHIC_AV_dout_nent(7),
      projin_7_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D4PHIC_enb,
      projin_7_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D4PHIC_V_readaddr,
      projin_7_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D4PHIC_V_dout,
      projin_7_mask_0_V                   => MPROJ_L1D1ABCD_D4PHIC_AV_dout_mask(0),
      projin_7_mask_1_V                   => MPROJ_L1D1ABCD_D4PHIC_AV_dout_mask(1),
      projin_7_nentries_0_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(0),
      projin_7_nentries_1_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(1),
      projin_7_nentries_2_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(2),
      projin_7_nentries_3_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(3),
      projin_7_nentries_4_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(4),
      projin_7_nentries_5_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(5),
      projin_7_nentries_6_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(6),
      projin_7_nentries_7_V               => MPROJ_L1D1ABCD_D4PHIC_AV_dout_nent(7),
      projin_8_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D4PHIC_enb,
      projin_8_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHIC_V_readaddr,
      projin_8_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D4PHIC_V_dout,
      projin_8_mask_0_V                   => MPROJ_L1D1EFGH_D4PHIC_AV_dout_mask(0),
      projin_8_mask_1_V                   => MPROJ_L1D1EFGH_D4PHIC_AV_dout_mask(1),
      projin_8_nentries_0_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(0),
      projin_8_nentries_1_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(1),
      projin_8_nentries_2_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(2),
      projin_8_nentries_3_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(3),
      projin_8_nentries_4_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(4),
      projin_8_nentries_5_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(5),
      projin_8_nentries_6_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(6),
      projin_8_nentries_7_V               => MPROJ_L1D1EFGH_D4PHIC_AV_dout_nent(7),
      projin_9_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D4PHIC_enb,
      projin_9_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHIC_V_readaddr,
      projin_9_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D4PHIC_V_dout,
      projin_9_mask_0_V                   => MPROJ_L2D1ABCD_D4PHIC_AV_dout_mask(0),
      projin_9_mask_1_V                   => MPROJ_L2D1ABCD_D4PHIC_AV_dout_mask(1),
      projin_9_nentries_0_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(0),
      projin_9_nentries_1_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(1),
      projin_9_nentries_2_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(2),
      projin_9_nentries_3_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(3),
      projin_9_nentries_4_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(4),
      projin_9_nentries_5_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(5),
      projin_9_nentries_6_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(6),
      projin_9_nentries_7_V               => MPROJ_L2D1ABCD_D4PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D4PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D4PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D4PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D4PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D4PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D4PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D4PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D4PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D4PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D4PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D4PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D4PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D4PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D4PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D4PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D4PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D4PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D4PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D4PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D4PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D4PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D4PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_D4PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D4PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D4PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D4PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D4PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D4PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D4PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D4PHIC_din
  );

  LATCH_MP_D4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D4PHID_bx,
      start => MP_D4PHID_start
  );

  MP_D4PHID : entity work.MP_D4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D4PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D4PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_L1L2G_D4PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_L1L2G_D4PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_L1L2G_D4PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_L1L2G_D4PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_L1L2G_D4PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_L1L2G_D4PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_L1L2HI_D4PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_L1L2HI_D4PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_L1L2HI_D4PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_L1L2HI_D4PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_L1L2HI_D4PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_L1L2HI_D4PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1L2JKL_D4PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1L2JKL_D4PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1L2JKL_D4PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1L2JKL_D4PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1L2JKL_D4PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1L2JKL_D4PHID_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L2L3ABCD_D4PHID_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L2L3ABCD_D4PHID_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L2L3ABCD_D4PHID_V_dout,
      projin_3_mask_0_V                   => MPROJ_L2L3ABCD_D4PHID_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L2L3ABCD_D4PHID_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L2L3ABCD_D4PHID_AV_dout_nent(7),
      projin_4_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D4PHID_enb,
      projin_4_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D4PHID_V_readaddr,
      projin_4_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D4PHID_V_dout,
      projin_4_mask_0_V                   => MPROJ_D1D2ABCD_D4PHID_AV_dout_mask(0),
      projin_4_mask_1_V                   => MPROJ_D1D2ABCD_D4PHID_AV_dout_mask(1),
      projin_4_nentries_0_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(0),
      projin_4_nentries_1_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(1),
      projin_4_nentries_2_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(2),
      projin_4_nentries_3_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(3),
      projin_4_nentries_4_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(4),
      projin_4_nentries_5_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(5),
      projin_4_nentries_6_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(6),
      projin_4_nentries_7_V               => MPROJ_D1D2ABCD_D4PHID_AV_dout_nent(7),
      projin_5_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D4PHID_enb,
      projin_5_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D4PHID_V_readaddr,
      projin_5_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D4PHID_V_dout,
      projin_5_mask_0_V                   => MPROJ_L1D1EFGH_D4PHID_AV_dout_mask(0),
      projin_5_mask_1_V                   => MPROJ_L1D1EFGH_D4PHID_AV_dout_mask(1),
      projin_5_nentries_0_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(0),
      projin_5_nentries_1_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(1),
      projin_5_nentries_2_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(2),
      projin_5_nentries_3_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(3),
      projin_5_nentries_4_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(4),
      projin_5_nentries_5_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(5),
      projin_5_nentries_6_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(6),
      projin_5_nentries_7_V               => MPROJ_L1D1EFGH_D4PHID_AV_dout_nent(7),
      projin_6_dataarray_data_V_ce0       => MPROJ_L2D1ABCD_D4PHID_enb,
      projin_6_dataarray_data_V_address0  => MPROJ_L2D1ABCD_D4PHID_V_readaddr,
      projin_6_dataarray_data_V_q0        => MPROJ_L2D1ABCD_D4PHID_V_dout,
      projin_6_mask_0_V                   => MPROJ_L2D1ABCD_D4PHID_AV_dout_mask(0),
      projin_6_mask_1_V                   => MPROJ_L2D1ABCD_D4PHID_AV_dout_mask(1),
      projin_6_nentries_0_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(0),
      projin_6_nentries_1_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(1),
      projin_6_nentries_2_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(2),
      projin_6_nentries_3_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(3),
      projin_6_nentries_4_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(4),
      projin_6_nentries_5_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(5),
      projin_6_nentries_6_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(6),
      projin_6_nentries_7_V               => MPROJ_L2D1ABCD_D4PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D4PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D4PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D4PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D4PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D4PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D4PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D4PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D4PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D4PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D4PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D4PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D4PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D4PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D4PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D4PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D4PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D4PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D4PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D4PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D4PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D4PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D4PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_D4PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D4PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D4PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D4PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D4PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D4PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D4PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D4PHID_din
  );

  LATCH_MP_D5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D5PHIA_bx,
      start => MP_D5PHIA_start
  );

  MP_D5PHIA : entity work.MP_D5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D5PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D5PHIA_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D5PHIA_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIA_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D5PHIA_V_dout,
      projin_0_mask_0_V                   => MPROJ_D1D2ABCD_D5PHIA_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_D1D2ABCD_D5PHIA_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_D1D2ABCD_D5PHIA_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D5PHIA_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIA_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D5PHIA_V_dout,
      projin_1_mask_0_V                   => MPROJ_D3D4ABCD_D5PHIA_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_D3D4ABCD_D5PHIA_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_D3D4ABCD_D5PHIA_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D5PHIA_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIA_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D5PHIA_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1D1ABCD_D5PHIA_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1D1ABCD_D5PHIA_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1D1ABCD_D5PHIA_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D5PHIAn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D5PHIAn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D5PHIAn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D5PHIAn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D5PHIAn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D5PHIAn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D5PHIAn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D5PHIAn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D5PHIAn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D5PHIAn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D5PHIAn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D5PHIAn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D5PHIAn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D5PHIAn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D5PHIAn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D5PHIAn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D5PHIAn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D5PHIAn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D5PHIAn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D5PHIAn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D5PHIAn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D5PHIAn2_enb,
      allstub_dataarray_data_V_address0  => AS_D5PHIAn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D5PHIAn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D5PHIA_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D5PHIA_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D5PHIA_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D5PHIA_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D5PHIA_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D5PHIA_din
  );

  LATCH_MP_D5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D5PHIB_bx,
      start => MP_D5PHIB_start
  );

  MP_D5PHIB : entity work.MP_D5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D5PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D5PHIB_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D5PHIB_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIB_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D5PHIB_V_dout,
      projin_0_mask_0_V                   => MPROJ_D1D2ABCD_D5PHIB_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_D1D2ABCD_D5PHIB_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_D1D2ABCD_D5PHIB_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D5PHIB_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIB_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D5PHIB_V_dout,
      projin_1_mask_0_V                   => MPROJ_D3D4ABCD_D5PHIB_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_D3D4ABCD_D5PHIB_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_D3D4ABCD_D5PHIB_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D5PHIB_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIB_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D5PHIB_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1D1ABCD_D5PHIB_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1D1ABCD_D5PHIB_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1D1ABCD_D5PHIB_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D5PHIB_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHIB_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D5PHIB_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1D1EFGH_D5PHIB_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1D1EFGH_D5PHIB_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1D1EFGH_D5PHIB_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D5PHIBn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D5PHIBn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D5PHIBn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D5PHIBn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D5PHIBn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D5PHIBn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D5PHIBn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D5PHIBn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D5PHIBn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D5PHIBn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D5PHIBn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D5PHIBn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D5PHIBn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D5PHIBn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D5PHIBn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D5PHIBn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D5PHIBn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D5PHIBn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D5PHIBn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D5PHIBn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D5PHIBn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D5PHIBn2_enb,
      allstub_dataarray_data_V_address0  => AS_D5PHIBn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D5PHIBn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D5PHIB_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D5PHIB_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D5PHIB_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D5PHIB_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D5PHIB_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D5PHIB_din
  );

  LATCH_MP_D5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D5PHIC_bx,
      start => MP_D5PHIC_start
  );

  MP_D5PHIC : entity work.MP_D5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D5PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D5PHIC_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D5PHIC_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHIC_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D5PHIC_V_dout,
      projin_0_mask_0_V                   => MPROJ_D1D2ABCD_D5PHIC_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_D1D2ABCD_D5PHIC_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_D1D2ABCD_D5PHIC_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D5PHIC_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHIC_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D5PHIC_V_dout,
      projin_1_mask_0_V                   => MPROJ_D3D4ABCD_D5PHIC_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_D3D4ABCD_D5PHIC_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_D3D4ABCD_D5PHIC_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1D1ABCD_D5PHIC_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1D1ABCD_D5PHIC_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1D1ABCD_D5PHIC_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1D1ABCD_D5PHIC_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1D1ABCD_D5PHIC_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1D1ABCD_D5PHIC_AV_dout_nent(7),
      projin_3_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D5PHIC_enb,
      projin_3_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHIC_V_readaddr,
      projin_3_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D5PHIC_V_dout,
      projin_3_mask_0_V                   => MPROJ_L1D1EFGH_D5PHIC_AV_dout_mask(0),
      projin_3_mask_1_V                   => MPROJ_L1D1EFGH_D5PHIC_AV_dout_mask(1),
      projin_3_nentries_0_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(0),
      projin_3_nentries_1_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(1),
      projin_3_nentries_2_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(2),
      projin_3_nentries_3_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(3),
      projin_3_nentries_4_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(4),
      projin_3_nentries_5_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(5),
      projin_3_nentries_6_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(6),
      projin_3_nentries_7_V               => MPROJ_L1D1EFGH_D5PHIC_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D5PHICn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D5PHICn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D5PHICn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D5PHICn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D5PHICn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D5PHICn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D5PHICn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D5PHICn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D5PHICn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D5PHICn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D5PHICn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D5PHICn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D5PHICn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D5PHICn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D5PHICn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D5PHICn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D5PHICn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D5PHICn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D5PHICn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D5PHICn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D5PHICn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D5PHICn2_enb,
      allstub_dataarray_data_V_address0  => AS_D5PHICn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D5PHICn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D5PHIC_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D5PHIC_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D5PHIC_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D5PHIC_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D5PHIC_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D5PHIC_din
  );

  LATCH_MP_D5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => PC_done,
      bx_out => PC_bx_out,
      bx => MP_D5PHID_bx,
      start => MP_D5PHID_start
  );

  MP_D5PHID : entity work.MP_D5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => MP_D5PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => MP_D5PHID_bx,
      projin_0_dataarray_data_V_ce0       => MPROJ_D1D2ABCD_D5PHID_enb,
      projin_0_dataarray_data_V_address0  => MPROJ_D1D2ABCD_D5PHID_V_readaddr,
      projin_0_dataarray_data_V_q0        => MPROJ_D1D2ABCD_D5PHID_V_dout,
      projin_0_mask_0_V                   => MPROJ_D1D2ABCD_D5PHID_AV_dout_mask(0),
      projin_0_mask_1_V                   => MPROJ_D1D2ABCD_D5PHID_AV_dout_mask(1),
      projin_0_nentries_0_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(0),
      projin_0_nentries_1_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(1),
      projin_0_nentries_2_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(2),
      projin_0_nentries_3_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(3),
      projin_0_nentries_4_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(4),
      projin_0_nentries_5_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(5),
      projin_0_nentries_6_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(6),
      projin_0_nentries_7_V               => MPROJ_D1D2ABCD_D5PHID_AV_dout_nent(7),
      projin_1_dataarray_data_V_ce0       => MPROJ_D3D4ABCD_D5PHID_enb,
      projin_1_dataarray_data_V_address0  => MPROJ_D3D4ABCD_D5PHID_V_readaddr,
      projin_1_dataarray_data_V_q0        => MPROJ_D3D4ABCD_D5PHID_V_dout,
      projin_1_mask_0_V                   => MPROJ_D3D4ABCD_D5PHID_AV_dout_mask(0),
      projin_1_mask_1_V                   => MPROJ_D3D4ABCD_D5PHID_AV_dout_mask(1),
      projin_1_nentries_0_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(0),
      projin_1_nentries_1_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(1),
      projin_1_nentries_2_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(2),
      projin_1_nentries_3_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(3),
      projin_1_nentries_4_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(4),
      projin_1_nentries_5_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(5),
      projin_1_nentries_6_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(6),
      projin_1_nentries_7_V               => MPROJ_D3D4ABCD_D5PHID_AV_dout_nent(7),
      projin_2_dataarray_data_V_ce0       => MPROJ_L1D1EFGH_D5PHID_enb,
      projin_2_dataarray_data_V_address0  => MPROJ_L1D1EFGH_D5PHID_V_readaddr,
      projin_2_dataarray_data_V_q0        => MPROJ_L1D1EFGH_D5PHID_V_dout,
      projin_2_mask_0_V                   => MPROJ_L1D1EFGH_D5PHID_AV_dout_mask(0),
      projin_2_mask_1_V                   => MPROJ_L1D1EFGH_D5PHID_AV_dout_mask(1),
      projin_2_nentries_0_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(0),
      projin_2_nentries_1_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(1),
      projin_2_nentries_2_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(2),
      projin_2_nentries_3_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(3),
      projin_2_nentries_4_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(4),
      projin_2_nentries_5_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(5),
      projin_2_nentries_6_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(6),
      projin_2_nentries_7_V               => MPROJ_L1D1EFGH_D5PHID_AV_dout_nent(7),
      instubdata_dataarray_0_data_V_ce0       => VMSME_D5PHIDn2_A_enb(0),
      instubdata_dataarray_0_data_V_address0  => VMSME_D5PHIDn2_AV_readaddr(0),
      instubdata_dataarray_0_data_V_q0        => VMSME_D5PHIDn2_AV_dout(0),
      instubdata_dataarray_1_data_V_ce0       => VMSME_D5PHIDn2_A_enb(1),
      instubdata_dataarray_1_data_V_address0  => VMSME_D5PHIDn2_AV_readaddr(1),
      instubdata_dataarray_1_data_V_q0        => VMSME_D5PHIDn2_AV_dout(1),
      instubdata_dataarray_2_data_V_ce0       => VMSME_D5PHIDn2_A_enb(2),
      instubdata_dataarray_2_data_V_address0  => VMSME_D5PHIDn2_AV_readaddr(2),
      instubdata_dataarray_2_data_V_q0        => VMSME_D5PHIDn2_AV_dout(2),
      instubdata_dataarray_3_data_V_ce0       => VMSME_D5PHIDn2_A_enb(3),
      instubdata_dataarray_3_data_V_address0  => VMSME_D5PHIDn2_AV_readaddr(3),
      instubdata_dataarray_3_data_V_q0        => VMSME_D5PHIDn2_AV_dout(3),
      instubdata_nentries_V_ce0 => VMSME_D5PHIDn2_enb_nent,
      instubdata_nentries_V_address0 => VMSME_D5PHIDn2_V_addr_nent,
      instubdata_nentries_V_q0 => VMSME_D5PHIDn2_AV_dout_nent,
      instubdata_binmaskA_V_address0 => VMSME_D5PHIDn2_V_addr_binmaskA,
      instubdata_binmaskA_V_ce0 => VMSME_D5PHIDn2_enb_binmaskA,
      instubdata_binmaskA_V_q0 => VMSME_D5PHIDn2_V_binmaskA,
      instubdata_binmaskB_V_address0 => VMSME_D5PHIDn2_V_addr_binmaskB,
      instubdata_binmaskB_V_ce0 => VMSME_D5PHIDn2_enb_binmaskB,
      instubdata_binmaskB_V_q0 => VMSME_D5PHIDn2_V_binmaskB,
      allstub_dataarray_data_V_ce0       => AS_D5PHIDn2_enb,
      allstub_dataarray_data_V_address0  => AS_D5PHIDn2_V_readaddr,
      allstub_dataarray_data_V_q0        => AS_D5PHIDn2_V_dout,
      fullmatch_0_dataarray_data_V_ce0       => open,
      fullmatch_0_dataarray_data_V_we0       => FM_AAAA_D5PHID_wea,
      fullmatch_0_dataarray_data_V_address0  => FM_AAAA_D5PHID_writeaddr,
      fullmatch_0_dataarray_data_V_d0        => FM_AAAA_D5PHID_din,
      fullmatch_1_dataarray_data_V_ce0       => open,
      fullmatch_1_dataarray_data_V_we0       => FM_BBBB_D5PHID_wea,
      fullmatch_1_dataarray_data_V_address0  => FM_BBBB_D5PHID_writeaddr,
      fullmatch_1_dataarray_data_V_d0        => FM_BBBB_D5PHID_din
  );

  LATCH_TB_AAAA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => MP_done,
      bx_out => MP_bx_out,
      bx => TB_AAAA_bx,
      start => TB_AAAA_start
  );

  TB_AAAA : entity work.TB_AAAA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TB_AAAA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TB_done,
      bx_V          => TB_AAAA_bx,
      bx_o_V        => TB_bx_out,
      bx_o_V_ap_vld => TB_bx_out_vld,
      trackletParameters1_0_dataarray_data_V_ce0       => MPAR_L1L2F_enb,
      trackletParameters1_0_dataarray_data_V_address0  => MPAR_L1L2F_V_readaddr,
      trackletParameters1_0_dataarray_data_V_q0        => MPAR_L1L2F_V_dout,
      trackletParameters1_1_dataarray_data_V_ce0       => MPAR_L1L2G_enb,
      trackletParameters1_1_dataarray_data_V_address0  => MPAR_L1L2G_V_readaddr,
      trackletParameters1_1_dataarray_data_V_q0        => MPAR_L1L2G_V_dout,
      trackletParameters2_0_dataarray_data_V_ce0       => MPAR_L1L2DE_enb,
      trackletParameters2_0_dataarray_data_V_address0  => MPAR_L1L2DE_V_readaddr,
      trackletParameters2_0_dataarray_data_V_q0        => MPAR_L1L2DE_V_dout,
      trackletParameters2_1_dataarray_data_V_ce0       => MPAR_L1L2HI_enb,
      trackletParameters2_1_dataarray_data_V_address0  => MPAR_L1L2HI_V_readaddr,
      trackletParameters2_1_dataarray_data_V_q0        => MPAR_L1L2HI_V_dout,
      trackletParameters3_0_dataarray_data_V_ce0       => MPAR_L1L2ABC_enb,
      trackletParameters3_0_dataarray_data_V_address0  => MPAR_L1L2ABC_V_readaddr,
      trackletParameters3_0_dataarray_data_V_q0        => MPAR_L1L2ABC_V_dout,
      trackletParameters3_1_dataarray_data_V_ce0       => MPAR_L1L2JKL_enb,
      trackletParameters3_1_dataarray_data_V_address0  => MPAR_L1L2JKL_V_readaddr,
      trackletParameters3_1_dataarray_data_V_q0        => MPAR_L1L2JKL_V_dout,
      trackletParameters4_0_dataarray_data_V_ce0       => MPAR_L2L3ABCD_enb,
      trackletParameters4_0_dataarray_data_V_address0  => MPAR_L2L3ABCD_V_readaddr,
      trackletParameters4_0_dataarray_data_V_q0        => MPAR_L2L3ABCD_V_dout,
      trackletParameters4_1_dataarray_data_V_ce0       => MPAR_L5L6ABCD_enb,
      trackletParameters4_1_dataarray_data_V_address0  => MPAR_L5L6ABCD_V_readaddr,
      trackletParameters4_1_dataarray_data_V_q0        => MPAR_L5L6ABCD_V_dout,
      trackletParameters4_2_dataarray_data_V_ce0       => MPAR_L2D1ABCD_enb,
      trackletParameters4_2_dataarray_data_V_address0  => MPAR_L2D1ABCD_V_readaddr,
      trackletParameters4_2_dataarray_data_V_q0        => MPAR_L2D1ABCD_V_dout,
      barrelFullMatches_0_dataarray_data_V_ce0       => FM_AAAA_L1PHIA_enb,
      barrelFullMatches_0_dataarray_data_V_address0  => FM_AAAA_L1PHIA_V_readaddr,
      barrelFullMatches_0_dataarray_data_V_q0        => FM_AAAA_L1PHIA_V_dout,
      barrelFullMatches_0_nentries_0_V               => FM_AAAA_L1PHIA_AV_dout_nent(0),
      barrelFullMatches_0_nentries_1_V               => FM_AAAA_L1PHIA_AV_dout_nent(1),
      barrelFullMatches_1_dataarray_data_V_ce0       => FM_AAAA_L1PHIB_enb,
      barrelFullMatches_1_dataarray_data_V_address0  => FM_AAAA_L1PHIB_V_readaddr,
      barrelFullMatches_1_dataarray_data_V_q0        => FM_AAAA_L1PHIB_V_dout,
      barrelFullMatches_1_nentries_0_V               => FM_AAAA_L1PHIB_AV_dout_nent(0),
      barrelFullMatches_1_nentries_1_V               => FM_AAAA_L1PHIB_AV_dout_nent(1),
      barrelFullMatches_2_dataarray_data_V_ce0       => FM_AAAA_L1PHIC_enb,
      barrelFullMatches_2_dataarray_data_V_address0  => FM_AAAA_L1PHIC_V_readaddr,
      barrelFullMatches_2_dataarray_data_V_q0        => FM_AAAA_L1PHIC_V_dout,
      barrelFullMatches_2_nentries_0_V               => FM_AAAA_L1PHIC_AV_dout_nent(0),
      barrelFullMatches_2_nentries_1_V               => FM_AAAA_L1PHIC_AV_dout_nent(1),
      barrelFullMatches_3_dataarray_data_V_ce0       => FM_AAAA_L1PHID_enb,
      barrelFullMatches_3_dataarray_data_V_address0  => FM_AAAA_L1PHID_V_readaddr,
      barrelFullMatches_3_dataarray_data_V_q0        => FM_AAAA_L1PHID_V_dout,
      barrelFullMatches_3_nentries_0_V               => FM_AAAA_L1PHID_AV_dout_nent(0),
      barrelFullMatches_3_nentries_1_V               => FM_AAAA_L1PHID_AV_dout_nent(1),
      barrelFullMatches_4_dataarray_data_V_ce0       => FM_AAAA_L1PHIE_enb,
      barrelFullMatches_4_dataarray_data_V_address0  => FM_AAAA_L1PHIE_V_readaddr,
      barrelFullMatches_4_dataarray_data_V_q0        => FM_AAAA_L1PHIE_V_dout,
      barrelFullMatches_4_nentries_0_V               => FM_AAAA_L1PHIE_AV_dout_nent(0),
      barrelFullMatches_4_nentries_1_V               => FM_AAAA_L1PHIE_AV_dout_nent(1),
      barrelFullMatches_5_dataarray_data_V_ce0       => FM_AAAA_L1PHIF_enb,
      barrelFullMatches_5_dataarray_data_V_address0  => FM_AAAA_L1PHIF_V_readaddr,
      barrelFullMatches_5_dataarray_data_V_q0        => FM_AAAA_L1PHIF_V_dout,
      barrelFullMatches_5_nentries_0_V               => FM_AAAA_L1PHIF_AV_dout_nent(0),
      barrelFullMatches_5_nentries_1_V               => FM_AAAA_L1PHIF_AV_dout_nent(1),
      barrelFullMatches_6_dataarray_data_V_ce0       => FM_AAAA_L1PHIG_enb,
      barrelFullMatches_6_dataarray_data_V_address0  => FM_AAAA_L1PHIG_V_readaddr,
      barrelFullMatches_6_dataarray_data_V_q0        => FM_AAAA_L1PHIG_V_dout,
      barrelFullMatches_6_nentries_0_V               => FM_AAAA_L1PHIG_AV_dout_nent(0),
      barrelFullMatches_6_nentries_1_V               => FM_AAAA_L1PHIG_AV_dout_nent(1),
      barrelFullMatches_7_dataarray_data_V_ce0       => FM_AAAA_L1PHIH_enb,
      barrelFullMatches_7_dataarray_data_V_address0  => FM_AAAA_L1PHIH_V_readaddr,
      barrelFullMatches_7_dataarray_data_V_q0        => FM_AAAA_L1PHIH_V_dout,
      barrelFullMatches_7_nentries_0_V               => FM_AAAA_L1PHIH_AV_dout_nent(0),
      barrelFullMatches_7_nentries_1_V               => FM_AAAA_L1PHIH_AV_dout_nent(1),
      barrelFullMatches_8_dataarray_data_V_ce0       => FM_AAAA_L2PHIA_enb,
      barrelFullMatches_8_dataarray_data_V_address0  => FM_AAAA_L2PHIA_V_readaddr,
      barrelFullMatches_8_dataarray_data_V_q0        => FM_AAAA_L2PHIA_V_dout,
      barrelFullMatches_8_nentries_0_V               => FM_AAAA_L2PHIA_AV_dout_nent(0),
      barrelFullMatches_8_nentries_1_V               => FM_AAAA_L2PHIA_AV_dout_nent(1),
      barrelFullMatches_9_dataarray_data_V_ce0       => FM_AAAA_L2PHIB_enb,
      barrelFullMatches_9_dataarray_data_V_address0  => FM_AAAA_L2PHIB_V_readaddr,
      barrelFullMatches_9_dataarray_data_V_q0        => FM_AAAA_L2PHIB_V_dout,
      barrelFullMatches_9_nentries_0_V               => FM_AAAA_L2PHIB_AV_dout_nent(0),
      barrelFullMatches_9_nentries_1_V               => FM_AAAA_L2PHIB_AV_dout_nent(1),
      barrelFullMatches_10_dataarray_data_V_ce0       => FM_AAAA_L2PHIC_enb,
      barrelFullMatches_10_dataarray_data_V_address0  => FM_AAAA_L2PHIC_V_readaddr,
      barrelFullMatches_10_dataarray_data_V_q0        => FM_AAAA_L2PHIC_V_dout,
      barrelFullMatches_10_nentries_0_V               => FM_AAAA_L2PHIC_AV_dout_nent(0),
      barrelFullMatches_10_nentries_1_V               => FM_AAAA_L2PHIC_AV_dout_nent(1),
      barrelFullMatches_11_dataarray_data_V_ce0       => FM_AAAA_L2PHID_enb,
      barrelFullMatches_11_dataarray_data_V_address0  => FM_AAAA_L2PHID_V_readaddr,
      barrelFullMatches_11_dataarray_data_V_q0        => FM_AAAA_L2PHID_V_dout,
      barrelFullMatches_11_nentries_0_V               => FM_AAAA_L2PHID_AV_dout_nent(0),
      barrelFullMatches_11_nentries_1_V               => FM_AAAA_L2PHID_AV_dout_nent(1),
      barrelFullMatches_12_dataarray_data_V_ce0       => FM_AAAA_L3PHIA_enb,
      barrelFullMatches_12_dataarray_data_V_address0  => FM_AAAA_L3PHIA_V_readaddr,
      barrelFullMatches_12_dataarray_data_V_q0        => FM_AAAA_L3PHIA_V_dout,
      barrelFullMatches_12_nentries_0_V               => FM_AAAA_L3PHIA_AV_dout_nent(0),
      barrelFullMatches_12_nentries_1_V               => FM_AAAA_L3PHIA_AV_dout_nent(1),
      barrelFullMatches_13_dataarray_data_V_ce0       => FM_AAAA_L3PHIB_enb,
      barrelFullMatches_13_dataarray_data_V_address0  => FM_AAAA_L3PHIB_V_readaddr,
      barrelFullMatches_13_dataarray_data_V_q0        => FM_AAAA_L3PHIB_V_dout,
      barrelFullMatches_13_nentries_0_V               => FM_AAAA_L3PHIB_AV_dout_nent(0),
      barrelFullMatches_13_nentries_1_V               => FM_AAAA_L3PHIB_AV_dout_nent(1),
      barrelFullMatches_14_dataarray_data_V_ce0       => FM_AAAA_L3PHIC_enb,
      barrelFullMatches_14_dataarray_data_V_address0  => FM_AAAA_L3PHIC_V_readaddr,
      barrelFullMatches_14_dataarray_data_V_q0        => FM_AAAA_L3PHIC_V_dout,
      barrelFullMatches_14_nentries_0_V               => FM_AAAA_L3PHIC_AV_dout_nent(0),
      barrelFullMatches_14_nentries_1_V               => FM_AAAA_L3PHIC_AV_dout_nent(1),
      barrelFullMatches_15_dataarray_data_V_ce0       => FM_AAAA_L3PHID_enb,
      barrelFullMatches_15_dataarray_data_V_address0  => FM_AAAA_L3PHID_V_readaddr,
      barrelFullMatches_15_dataarray_data_V_q0        => FM_AAAA_L3PHID_V_dout,
      barrelFullMatches_15_nentries_0_V               => FM_AAAA_L3PHID_AV_dout_nent(0),
      barrelFullMatches_15_nentries_1_V               => FM_AAAA_L3PHID_AV_dout_nent(1),
      barrelFullMatches_16_dataarray_data_V_ce0       => FM_AAAA_L4PHIA_enb,
      barrelFullMatches_16_dataarray_data_V_address0  => FM_AAAA_L4PHIA_V_readaddr,
      barrelFullMatches_16_dataarray_data_V_q0        => FM_AAAA_L4PHIA_V_dout,
      barrelFullMatches_16_nentries_0_V               => FM_AAAA_L4PHIA_AV_dout_nent(0),
      barrelFullMatches_16_nentries_1_V               => FM_AAAA_L4PHIA_AV_dout_nent(1),
      barrelFullMatches_17_dataarray_data_V_ce0       => FM_AAAA_L4PHIB_enb,
      barrelFullMatches_17_dataarray_data_V_address0  => FM_AAAA_L4PHIB_V_readaddr,
      barrelFullMatches_17_dataarray_data_V_q0        => FM_AAAA_L4PHIB_V_dout,
      barrelFullMatches_17_nentries_0_V               => FM_AAAA_L4PHIB_AV_dout_nent(0),
      barrelFullMatches_17_nentries_1_V               => FM_AAAA_L4PHIB_AV_dout_nent(1),
      barrelFullMatches_18_dataarray_data_V_ce0       => FM_AAAA_L4PHIC_enb,
      barrelFullMatches_18_dataarray_data_V_address0  => FM_AAAA_L4PHIC_V_readaddr,
      barrelFullMatches_18_dataarray_data_V_q0        => FM_AAAA_L4PHIC_V_dout,
      barrelFullMatches_18_nentries_0_V               => FM_AAAA_L4PHIC_AV_dout_nent(0),
      barrelFullMatches_18_nentries_1_V               => FM_AAAA_L4PHIC_AV_dout_nent(1),
      barrelFullMatches_19_dataarray_data_V_ce0       => FM_AAAA_L4PHID_enb,
      barrelFullMatches_19_dataarray_data_V_address0  => FM_AAAA_L4PHID_V_readaddr,
      barrelFullMatches_19_dataarray_data_V_q0        => FM_AAAA_L4PHID_V_dout,
      barrelFullMatches_19_nentries_0_V               => FM_AAAA_L4PHID_AV_dout_nent(0),
      barrelFullMatches_19_nentries_1_V               => FM_AAAA_L4PHID_AV_dout_nent(1),
      barrelFullMatches_20_dataarray_data_V_ce0       => FM_AAAA_L5PHIA_enb,
      barrelFullMatches_20_dataarray_data_V_address0  => FM_AAAA_L5PHIA_V_readaddr,
      barrelFullMatches_20_dataarray_data_V_q0        => FM_AAAA_L5PHIA_V_dout,
      barrelFullMatches_20_nentries_0_V               => FM_AAAA_L5PHIA_AV_dout_nent(0),
      barrelFullMatches_20_nentries_1_V               => FM_AAAA_L5PHIA_AV_dout_nent(1),
      barrelFullMatches_21_dataarray_data_V_ce0       => FM_AAAA_L5PHIB_enb,
      barrelFullMatches_21_dataarray_data_V_address0  => FM_AAAA_L5PHIB_V_readaddr,
      barrelFullMatches_21_dataarray_data_V_q0        => FM_AAAA_L5PHIB_V_dout,
      barrelFullMatches_21_nentries_0_V               => FM_AAAA_L5PHIB_AV_dout_nent(0),
      barrelFullMatches_21_nentries_1_V               => FM_AAAA_L5PHIB_AV_dout_nent(1),
      barrelFullMatches_22_dataarray_data_V_ce0       => FM_AAAA_L5PHIC_enb,
      barrelFullMatches_22_dataarray_data_V_address0  => FM_AAAA_L5PHIC_V_readaddr,
      barrelFullMatches_22_dataarray_data_V_q0        => FM_AAAA_L5PHIC_V_dout,
      barrelFullMatches_22_nentries_0_V               => FM_AAAA_L5PHIC_AV_dout_nent(0),
      barrelFullMatches_22_nentries_1_V               => FM_AAAA_L5PHIC_AV_dout_nent(1),
      barrelFullMatches_23_dataarray_data_V_ce0       => FM_AAAA_L5PHID_enb,
      barrelFullMatches_23_dataarray_data_V_address0  => FM_AAAA_L5PHID_V_readaddr,
      barrelFullMatches_23_dataarray_data_V_q0        => FM_AAAA_L5PHID_V_dout,
      barrelFullMatches_23_nentries_0_V               => FM_AAAA_L5PHID_AV_dout_nent(0),
      barrelFullMatches_23_nentries_1_V               => FM_AAAA_L5PHID_AV_dout_nent(1),
      barrelFullMatches_24_dataarray_data_V_ce0       => FM_AAAA_L6PHIA_enb,
      barrelFullMatches_24_dataarray_data_V_address0  => FM_AAAA_L6PHIA_V_readaddr,
      barrelFullMatches_24_dataarray_data_V_q0        => FM_AAAA_L6PHIA_V_dout,
      barrelFullMatches_24_nentries_0_V               => FM_AAAA_L6PHIA_AV_dout_nent(0),
      barrelFullMatches_24_nentries_1_V               => FM_AAAA_L6PHIA_AV_dout_nent(1),
      barrelFullMatches_25_dataarray_data_V_ce0       => FM_AAAA_L6PHIB_enb,
      barrelFullMatches_25_dataarray_data_V_address0  => FM_AAAA_L6PHIB_V_readaddr,
      barrelFullMatches_25_dataarray_data_V_q0        => FM_AAAA_L6PHIB_V_dout,
      barrelFullMatches_25_nentries_0_V               => FM_AAAA_L6PHIB_AV_dout_nent(0),
      barrelFullMatches_25_nentries_1_V               => FM_AAAA_L6PHIB_AV_dout_nent(1),
      barrelFullMatches_26_dataarray_data_V_ce0       => FM_AAAA_L6PHIC_enb,
      barrelFullMatches_26_dataarray_data_V_address0  => FM_AAAA_L6PHIC_V_readaddr,
      barrelFullMatches_26_dataarray_data_V_q0        => FM_AAAA_L6PHIC_V_dout,
      barrelFullMatches_26_nentries_0_V               => FM_AAAA_L6PHIC_AV_dout_nent(0),
      barrelFullMatches_26_nentries_1_V               => FM_AAAA_L6PHIC_AV_dout_nent(1),
      barrelFullMatches_27_dataarray_data_V_ce0       => FM_AAAA_L6PHID_enb,
      barrelFullMatches_27_dataarray_data_V_address0  => FM_AAAA_L6PHID_V_readaddr,
      barrelFullMatches_27_dataarray_data_V_q0        => FM_AAAA_L6PHID_V_dout,
      barrelFullMatches_27_nentries_0_V               => FM_AAAA_L6PHID_AV_dout_nent(0),
      barrelFullMatches_27_nentries_1_V               => FM_AAAA_L6PHID_AV_dout_nent(1),
      diskFullMatches_0_dataarray_data_V_ce0       => FM_AAAA_D1PHIA_enb,
      diskFullMatches_0_dataarray_data_V_address0  => FM_AAAA_D1PHIA_V_readaddr,
      diskFullMatches_0_dataarray_data_V_q0        => FM_AAAA_D1PHIA_V_dout,
      diskFullMatches_0_nentries_0_V               => FM_AAAA_D1PHIA_AV_dout_nent(0),
      diskFullMatches_0_nentries_1_V               => FM_AAAA_D1PHIA_AV_dout_nent(1),
      diskFullMatches_1_dataarray_data_V_ce0       => FM_AAAA_D1PHIB_enb,
      diskFullMatches_1_dataarray_data_V_address0  => FM_AAAA_D1PHIB_V_readaddr,
      diskFullMatches_1_dataarray_data_V_q0        => FM_AAAA_D1PHIB_V_dout,
      diskFullMatches_1_nentries_0_V               => FM_AAAA_D1PHIB_AV_dout_nent(0),
      diskFullMatches_1_nentries_1_V               => FM_AAAA_D1PHIB_AV_dout_nent(1),
      diskFullMatches_2_dataarray_data_V_ce0       => FM_AAAA_D1PHIC_enb,
      diskFullMatches_2_dataarray_data_V_address0  => FM_AAAA_D1PHIC_V_readaddr,
      diskFullMatches_2_dataarray_data_V_q0        => FM_AAAA_D1PHIC_V_dout,
      diskFullMatches_2_nentries_0_V               => FM_AAAA_D1PHIC_AV_dout_nent(0),
      diskFullMatches_2_nentries_1_V               => FM_AAAA_D1PHIC_AV_dout_nent(1),
      diskFullMatches_3_dataarray_data_V_ce0       => FM_AAAA_D1PHID_enb,
      diskFullMatches_3_dataarray_data_V_address0  => FM_AAAA_D1PHID_V_readaddr,
      diskFullMatches_3_dataarray_data_V_q0        => FM_AAAA_D1PHID_V_dout,
      diskFullMatches_3_nentries_0_V               => FM_AAAA_D1PHID_AV_dout_nent(0),
      diskFullMatches_3_nentries_1_V               => FM_AAAA_D1PHID_AV_dout_nent(1),
      diskFullMatches_4_dataarray_data_V_ce0       => FM_AAAA_D2PHIA_enb,
      diskFullMatches_4_dataarray_data_V_address0  => FM_AAAA_D2PHIA_V_readaddr,
      diskFullMatches_4_dataarray_data_V_q0        => FM_AAAA_D2PHIA_V_dout,
      diskFullMatches_4_nentries_0_V               => FM_AAAA_D2PHIA_AV_dout_nent(0),
      diskFullMatches_4_nentries_1_V               => FM_AAAA_D2PHIA_AV_dout_nent(1),
      diskFullMatches_5_dataarray_data_V_ce0       => FM_AAAA_D2PHIB_enb,
      diskFullMatches_5_dataarray_data_V_address0  => FM_AAAA_D2PHIB_V_readaddr,
      diskFullMatches_5_dataarray_data_V_q0        => FM_AAAA_D2PHIB_V_dout,
      diskFullMatches_5_nentries_0_V               => FM_AAAA_D2PHIB_AV_dout_nent(0),
      diskFullMatches_5_nentries_1_V               => FM_AAAA_D2PHIB_AV_dout_nent(1),
      diskFullMatches_6_dataarray_data_V_ce0       => FM_AAAA_D2PHIC_enb,
      diskFullMatches_6_dataarray_data_V_address0  => FM_AAAA_D2PHIC_V_readaddr,
      diskFullMatches_6_dataarray_data_V_q0        => FM_AAAA_D2PHIC_V_dout,
      diskFullMatches_6_nentries_0_V               => FM_AAAA_D2PHIC_AV_dout_nent(0),
      diskFullMatches_6_nentries_1_V               => FM_AAAA_D2PHIC_AV_dout_nent(1),
      diskFullMatches_7_dataarray_data_V_ce0       => FM_AAAA_D2PHID_enb,
      diskFullMatches_7_dataarray_data_V_address0  => FM_AAAA_D2PHID_V_readaddr,
      diskFullMatches_7_dataarray_data_V_q0        => FM_AAAA_D2PHID_V_dout,
      diskFullMatches_7_nentries_0_V               => FM_AAAA_D2PHID_AV_dout_nent(0),
      diskFullMatches_7_nentries_1_V               => FM_AAAA_D2PHID_AV_dout_nent(1),
      diskFullMatches_8_dataarray_data_V_ce0       => FM_AAAA_D3PHIA_enb,
      diskFullMatches_8_dataarray_data_V_address0  => FM_AAAA_D3PHIA_V_readaddr,
      diskFullMatches_8_dataarray_data_V_q0        => FM_AAAA_D3PHIA_V_dout,
      diskFullMatches_8_nentries_0_V               => FM_AAAA_D3PHIA_AV_dout_nent(0),
      diskFullMatches_8_nentries_1_V               => FM_AAAA_D3PHIA_AV_dout_nent(1),
      diskFullMatches_9_dataarray_data_V_ce0       => FM_AAAA_D3PHIB_enb,
      diskFullMatches_9_dataarray_data_V_address0  => FM_AAAA_D3PHIB_V_readaddr,
      diskFullMatches_9_dataarray_data_V_q0        => FM_AAAA_D3PHIB_V_dout,
      diskFullMatches_9_nentries_0_V               => FM_AAAA_D3PHIB_AV_dout_nent(0),
      diskFullMatches_9_nentries_1_V               => FM_AAAA_D3PHIB_AV_dout_nent(1),
      diskFullMatches_10_dataarray_data_V_ce0       => FM_AAAA_D3PHIC_enb,
      diskFullMatches_10_dataarray_data_V_address0  => FM_AAAA_D3PHIC_V_readaddr,
      diskFullMatches_10_dataarray_data_V_q0        => FM_AAAA_D3PHIC_V_dout,
      diskFullMatches_10_nentries_0_V               => FM_AAAA_D3PHIC_AV_dout_nent(0),
      diskFullMatches_10_nentries_1_V               => FM_AAAA_D3PHIC_AV_dout_nent(1),
      diskFullMatches_11_dataarray_data_V_ce0       => FM_AAAA_D3PHID_enb,
      diskFullMatches_11_dataarray_data_V_address0  => FM_AAAA_D3PHID_V_readaddr,
      diskFullMatches_11_dataarray_data_V_q0        => FM_AAAA_D3PHID_V_dout,
      diskFullMatches_11_nentries_0_V               => FM_AAAA_D3PHID_AV_dout_nent(0),
      diskFullMatches_11_nentries_1_V               => FM_AAAA_D3PHID_AV_dout_nent(1),
      diskFullMatches_12_dataarray_data_V_ce0       => FM_AAAA_D4PHIA_enb,
      diskFullMatches_12_dataarray_data_V_address0  => FM_AAAA_D4PHIA_V_readaddr,
      diskFullMatches_12_dataarray_data_V_q0        => FM_AAAA_D4PHIA_V_dout,
      diskFullMatches_12_nentries_0_V               => FM_AAAA_D4PHIA_AV_dout_nent(0),
      diskFullMatches_12_nentries_1_V               => FM_AAAA_D4PHIA_AV_dout_nent(1),
      diskFullMatches_13_dataarray_data_V_ce0       => FM_AAAA_D4PHIB_enb,
      diskFullMatches_13_dataarray_data_V_address0  => FM_AAAA_D4PHIB_V_readaddr,
      diskFullMatches_13_dataarray_data_V_q0        => FM_AAAA_D4PHIB_V_dout,
      diskFullMatches_13_nentries_0_V               => FM_AAAA_D4PHIB_AV_dout_nent(0),
      diskFullMatches_13_nentries_1_V               => FM_AAAA_D4PHIB_AV_dout_nent(1),
      diskFullMatches_14_dataarray_data_V_ce0       => FM_AAAA_D4PHIC_enb,
      diskFullMatches_14_dataarray_data_V_address0  => FM_AAAA_D4PHIC_V_readaddr,
      diskFullMatches_14_dataarray_data_V_q0        => FM_AAAA_D4PHIC_V_dout,
      diskFullMatches_14_nentries_0_V               => FM_AAAA_D4PHIC_AV_dout_nent(0),
      diskFullMatches_14_nentries_1_V               => FM_AAAA_D4PHIC_AV_dout_nent(1),
      diskFullMatches_15_dataarray_data_V_ce0       => FM_AAAA_D4PHID_enb,
      diskFullMatches_15_dataarray_data_V_address0  => FM_AAAA_D4PHID_V_readaddr,
      diskFullMatches_15_dataarray_data_V_q0        => FM_AAAA_D4PHID_V_dout,
      diskFullMatches_15_nentries_0_V               => FM_AAAA_D4PHID_AV_dout_nent(0),
      diskFullMatches_15_nentries_1_V               => FM_AAAA_D4PHID_AV_dout_nent(1),
      diskFullMatches_16_dataarray_data_V_ce0       => FM_AAAA_D5PHIA_enb,
      diskFullMatches_16_dataarray_data_V_address0  => FM_AAAA_D5PHIA_V_readaddr,
      diskFullMatches_16_dataarray_data_V_q0        => FM_AAAA_D5PHIA_V_dout,
      diskFullMatches_16_nentries_0_V               => FM_AAAA_D5PHIA_AV_dout_nent(0),
      diskFullMatches_16_nentries_1_V               => FM_AAAA_D5PHIA_AV_dout_nent(1),
      diskFullMatches_17_dataarray_data_V_ce0       => FM_AAAA_D5PHIB_enb,
      diskFullMatches_17_dataarray_data_V_address0  => FM_AAAA_D5PHIB_V_readaddr,
      diskFullMatches_17_dataarray_data_V_q0        => FM_AAAA_D5PHIB_V_dout,
      diskFullMatches_17_nentries_0_V               => FM_AAAA_D5PHIB_AV_dout_nent(0),
      diskFullMatches_17_nentries_1_V               => FM_AAAA_D5PHIB_AV_dout_nent(1),
      diskFullMatches_18_dataarray_data_V_ce0       => FM_AAAA_D5PHIC_enb,
      diskFullMatches_18_dataarray_data_V_address0  => FM_AAAA_D5PHIC_V_readaddr,
      diskFullMatches_18_dataarray_data_V_q0        => FM_AAAA_D5PHIC_V_dout,
      diskFullMatches_18_nentries_0_V               => FM_AAAA_D5PHIC_AV_dout_nent(0),
      diskFullMatches_18_nentries_1_V               => FM_AAAA_D5PHIC_AV_dout_nent(1),
      diskFullMatches_19_dataarray_data_V_ce0       => FM_AAAA_D5PHID_enb,
      diskFullMatches_19_dataarray_data_V_address0  => FM_AAAA_D5PHID_V_readaddr,
      diskFullMatches_19_dataarray_data_V_q0        => FM_AAAA_D5PHID_V_dout,
      diskFullMatches_19_nentries_0_V               => FM_AAAA_D5PHID_AV_dout_nent(0),
      diskFullMatches_19_nentries_1_V               => FM_AAAA_D5PHID_AV_dout_nent(1),
      trackWord_V_din       => TW_AAAA_stream_AV_din,
      trackWord_V_full_n    => TW_AAAA_stream_A_full_neg,
      trackWord_V_write     => TW_AAAA_stream_A_write,
      barrelStubWords_0_V_din       => BW_AAAA_L1_stream_AV_din,
      barrelStubWords_0_V_full_n    => BW_AAAA_L1_stream_A_full_neg,
      barrelStubWords_0_V_write     => BW_AAAA_L1_stream_A_write,
      barrelStubWords_1_V_din       => BW_AAAA_L2_stream_AV_din,
      barrelStubWords_1_V_full_n    => BW_AAAA_L2_stream_A_full_neg,
      barrelStubWords_1_V_write     => BW_AAAA_L2_stream_A_write,
      barrelStubWords_2_V_din       => BW_AAAA_L3_stream_AV_din,
      barrelStubWords_2_V_full_n    => BW_AAAA_L3_stream_A_full_neg,
      barrelStubWords_2_V_write     => BW_AAAA_L3_stream_A_write,
      barrelStubWords_3_V_din       => BW_AAAA_L4_stream_AV_din,
      barrelStubWords_3_V_full_n    => BW_AAAA_L4_stream_A_full_neg,
      barrelStubWords_3_V_write     => BW_AAAA_L4_stream_A_write,
      barrelStubWords_4_V_din       => BW_AAAA_L5_stream_AV_din,
      barrelStubWords_4_V_full_n    => BW_AAAA_L5_stream_A_full_neg,
      barrelStubWords_4_V_write     => BW_AAAA_L5_stream_A_write,
      barrelStubWords_5_V_din       => BW_AAAA_L6_stream_AV_din,
      barrelStubWords_5_V_full_n    => BW_AAAA_L6_stream_A_full_neg,
      barrelStubWords_5_V_write     => BW_AAAA_L6_stream_A_write,
      diskStubWords_0_V_din       => DW_AAAA_D1_stream_AV_din,
      diskStubWords_0_V_full_n    => DW_AAAA_D1_stream_A_full_neg,
      diskStubWords_0_V_write     => DW_AAAA_D1_stream_A_write,
      diskStubWords_1_V_din       => DW_AAAA_D2_stream_AV_din,
      diskStubWords_1_V_full_n    => DW_AAAA_D2_stream_A_full_neg,
      diskStubWords_1_V_write     => DW_AAAA_D2_stream_A_write,
      diskStubWords_2_V_din       => DW_AAAA_D3_stream_AV_din,
      diskStubWords_2_V_full_n    => DW_AAAA_D3_stream_A_full_neg,
      diskStubWords_2_V_write     => DW_AAAA_D3_stream_A_write,
      diskStubWords_3_V_din       => DW_AAAA_D4_stream_AV_din,
      diskStubWords_3_V_full_n    => DW_AAAA_D4_stream_A_full_neg,
      diskStubWords_3_V_write     => DW_AAAA_D4_stream_A_write,
      diskStubWords_4_V_din       => DW_AAAA_D5_stream_AV_din,
      diskStubWords_4_V_full_n    => DW_AAAA_D5_stream_A_full_neg,
      diskStubWords_4_V_write     => DW_AAAA_D5_stream_A_write,
      done        => TB_AAAA_last_track,
      done_ap_vld => TB_AAAA_last_track_vld
  );

  LATCH_TB_BBBB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => MP_done,
      bx_out => MP_bx_out,
      bx => TB_BBBB_bx,
      start => TB_BBBB_start
  );

  TB_BBBB : entity work.TB_BBBB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TB_BBBB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TB_BBBB_bx,
      trackletParameters2_0_dataarray_data_V_ce0       => MPAR_L3L4AB_enb,
      trackletParameters2_0_dataarray_data_V_address0  => MPAR_L3L4AB_V_readaddr,
      trackletParameters2_0_dataarray_data_V_q0        => MPAR_L3L4AB_V_dout,
      trackletParameters2_1_dataarray_data_V_ce0       => MPAR_L3L4CD_enb,
      trackletParameters2_1_dataarray_data_V_address0  => MPAR_L3L4CD_V_readaddr,
      trackletParameters2_1_dataarray_data_V_q0        => MPAR_L3L4CD_V_dout,
      trackletParameters4_0_dataarray_data_V_ce0       => MPAR_D1D2ABCD_enb,
      trackletParameters4_0_dataarray_data_V_address0  => MPAR_D1D2ABCD_V_readaddr,
      trackletParameters4_0_dataarray_data_V_q0        => MPAR_D1D2ABCD_V_dout,
      trackletParameters4_1_dataarray_data_V_ce0       => MPAR_D3D4ABCD_enb,
      trackletParameters4_1_dataarray_data_V_address0  => MPAR_D3D4ABCD_V_readaddr,
      trackletParameters4_1_dataarray_data_V_q0        => MPAR_D3D4ABCD_V_dout,
      trackletParameters4_2_dataarray_data_V_ce0       => MPAR_L1D1ABCD_enb,
      trackletParameters4_2_dataarray_data_V_address0  => MPAR_L1D1ABCD_V_readaddr,
      trackletParameters4_2_dataarray_data_V_q0        => MPAR_L1D1ABCD_V_dout,
      trackletParameters4_3_dataarray_data_V_ce0       => MPAR_L1D1EFGH_enb,
      trackletParameters4_3_dataarray_data_V_address0  => MPAR_L1D1EFGH_V_readaddr,
      trackletParameters4_3_dataarray_data_V_q0        => MPAR_L1D1EFGH_V_dout,
      barrelFullMatches_0_dataarray_data_V_ce0       => FM_BBBB_L1PHIA_enb,
      barrelFullMatches_0_dataarray_data_V_address0  => FM_BBBB_L1PHIA_V_readaddr,
      barrelFullMatches_0_dataarray_data_V_q0        => FM_BBBB_L1PHIA_V_dout,
      barrelFullMatches_0_nentries_0_V               => FM_BBBB_L1PHIA_AV_dout_nent(0),
      barrelFullMatches_0_nentries_1_V               => FM_BBBB_L1PHIA_AV_dout_nent(1),
      barrelFullMatches_1_dataarray_data_V_ce0       => FM_BBBB_L1PHIB_enb,
      barrelFullMatches_1_dataarray_data_V_address0  => FM_BBBB_L1PHIB_V_readaddr,
      barrelFullMatches_1_dataarray_data_V_q0        => FM_BBBB_L1PHIB_V_dout,
      barrelFullMatches_1_nentries_0_V               => FM_BBBB_L1PHIB_AV_dout_nent(0),
      barrelFullMatches_1_nentries_1_V               => FM_BBBB_L1PHIB_AV_dout_nent(1),
      barrelFullMatches_2_dataarray_data_V_ce0       => FM_BBBB_L1PHIC_enb,
      barrelFullMatches_2_dataarray_data_V_address0  => FM_BBBB_L1PHIC_V_readaddr,
      barrelFullMatches_2_dataarray_data_V_q0        => FM_BBBB_L1PHIC_V_dout,
      barrelFullMatches_2_nentries_0_V               => FM_BBBB_L1PHIC_AV_dout_nent(0),
      barrelFullMatches_2_nentries_1_V               => FM_BBBB_L1PHIC_AV_dout_nent(1),
      barrelFullMatches_3_dataarray_data_V_ce0       => FM_BBBB_L1PHID_enb,
      barrelFullMatches_3_dataarray_data_V_address0  => FM_BBBB_L1PHID_V_readaddr,
      barrelFullMatches_3_dataarray_data_V_q0        => FM_BBBB_L1PHID_V_dout,
      barrelFullMatches_3_nentries_0_V               => FM_BBBB_L1PHID_AV_dout_nent(0),
      barrelFullMatches_3_nentries_1_V               => FM_BBBB_L1PHID_AV_dout_nent(1),
      barrelFullMatches_4_dataarray_data_V_ce0       => FM_BBBB_L1PHIE_enb,
      barrelFullMatches_4_dataarray_data_V_address0  => FM_BBBB_L1PHIE_V_readaddr,
      barrelFullMatches_4_dataarray_data_V_q0        => FM_BBBB_L1PHIE_V_dout,
      barrelFullMatches_4_nentries_0_V               => FM_BBBB_L1PHIE_AV_dout_nent(0),
      barrelFullMatches_4_nentries_1_V               => FM_BBBB_L1PHIE_AV_dout_nent(1),
      barrelFullMatches_5_dataarray_data_V_ce0       => FM_BBBB_L1PHIF_enb,
      barrelFullMatches_5_dataarray_data_V_address0  => FM_BBBB_L1PHIF_V_readaddr,
      barrelFullMatches_5_dataarray_data_V_q0        => FM_BBBB_L1PHIF_V_dout,
      barrelFullMatches_5_nentries_0_V               => FM_BBBB_L1PHIF_AV_dout_nent(0),
      barrelFullMatches_5_nentries_1_V               => FM_BBBB_L1PHIF_AV_dout_nent(1),
      barrelFullMatches_6_dataarray_data_V_ce0       => FM_BBBB_L1PHIG_enb,
      barrelFullMatches_6_dataarray_data_V_address0  => FM_BBBB_L1PHIG_V_readaddr,
      barrelFullMatches_6_dataarray_data_V_q0        => FM_BBBB_L1PHIG_V_dout,
      barrelFullMatches_6_nentries_0_V               => FM_BBBB_L1PHIG_AV_dout_nent(0),
      barrelFullMatches_6_nentries_1_V               => FM_BBBB_L1PHIG_AV_dout_nent(1),
      barrelFullMatches_7_dataarray_data_V_ce0       => FM_BBBB_L1PHIH_enb,
      barrelFullMatches_7_dataarray_data_V_address0  => FM_BBBB_L1PHIH_V_readaddr,
      barrelFullMatches_7_dataarray_data_V_q0        => FM_BBBB_L1PHIH_V_dout,
      barrelFullMatches_7_nentries_0_V               => FM_BBBB_L1PHIH_AV_dout_nent(0),
      barrelFullMatches_7_nentries_1_V               => FM_BBBB_L1PHIH_AV_dout_nent(1),
      barrelFullMatches_8_dataarray_data_V_ce0       => FM_BBBB_L2PHIA_enb,
      barrelFullMatches_8_dataarray_data_V_address0  => FM_BBBB_L2PHIA_V_readaddr,
      barrelFullMatches_8_dataarray_data_V_q0        => FM_BBBB_L2PHIA_V_dout,
      barrelFullMatches_8_nentries_0_V               => FM_BBBB_L2PHIA_AV_dout_nent(0),
      barrelFullMatches_8_nentries_1_V               => FM_BBBB_L2PHIA_AV_dout_nent(1),
      barrelFullMatches_9_dataarray_data_V_ce0       => FM_BBBB_L2PHIB_enb,
      barrelFullMatches_9_dataarray_data_V_address0  => FM_BBBB_L2PHIB_V_readaddr,
      barrelFullMatches_9_dataarray_data_V_q0        => FM_BBBB_L2PHIB_V_dout,
      barrelFullMatches_9_nentries_0_V               => FM_BBBB_L2PHIB_AV_dout_nent(0),
      barrelFullMatches_9_nentries_1_V               => FM_BBBB_L2PHIB_AV_dout_nent(1),
      barrelFullMatches_10_dataarray_data_V_ce0       => FM_BBBB_L2PHIC_enb,
      barrelFullMatches_10_dataarray_data_V_address0  => FM_BBBB_L2PHIC_V_readaddr,
      barrelFullMatches_10_dataarray_data_V_q0        => FM_BBBB_L2PHIC_V_dout,
      barrelFullMatches_10_nentries_0_V               => FM_BBBB_L2PHIC_AV_dout_nent(0),
      barrelFullMatches_10_nentries_1_V               => FM_BBBB_L2PHIC_AV_dout_nent(1),
      barrelFullMatches_11_dataarray_data_V_ce0       => FM_BBBB_L2PHID_enb,
      barrelFullMatches_11_dataarray_data_V_address0  => FM_BBBB_L2PHID_V_readaddr,
      barrelFullMatches_11_dataarray_data_V_q0        => FM_BBBB_L2PHID_V_dout,
      barrelFullMatches_11_nentries_0_V               => FM_BBBB_L2PHID_AV_dout_nent(0),
      barrelFullMatches_11_nentries_1_V               => FM_BBBB_L2PHID_AV_dout_nent(1),
      barrelFullMatches_12_dataarray_data_V_ce0       => FM_BBBB_L3PHIA_enb,
      barrelFullMatches_12_dataarray_data_V_address0  => FM_BBBB_L3PHIA_V_readaddr,
      barrelFullMatches_12_dataarray_data_V_q0        => FM_BBBB_L3PHIA_V_dout,
      barrelFullMatches_12_nentries_0_V               => FM_BBBB_L3PHIA_AV_dout_nent(0),
      barrelFullMatches_12_nentries_1_V               => FM_BBBB_L3PHIA_AV_dout_nent(1),
      barrelFullMatches_13_dataarray_data_V_ce0       => FM_BBBB_L3PHIB_enb,
      barrelFullMatches_13_dataarray_data_V_address0  => FM_BBBB_L3PHIB_V_readaddr,
      barrelFullMatches_13_dataarray_data_V_q0        => FM_BBBB_L3PHIB_V_dout,
      barrelFullMatches_13_nentries_0_V               => FM_BBBB_L3PHIB_AV_dout_nent(0),
      barrelFullMatches_13_nentries_1_V               => FM_BBBB_L3PHIB_AV_dout_nent(1),
      barrelFullMatches_14_dataarray_data_V_ce0       => FM_BBBB_L3PHIC_enb,
      barrelFullMatches_14_dataarray_data_V_address0  => FM_BBBB_L3PHIC_V_readaddr,
      barrelFullMatches_14_dataarray_data_V_q0        => FM_BBBB_L3PHIC_V_dout,
      barrelFullMatches_14_nentries_0_V               => FM_BBBB_L3PHIC_AV_dout_nent(0),
      barrelFullMatches_14_nentries_1_V               => FM_BBBB_L3PHIC_AV_dout_nent(1),
      barrelFullMatches_15_dataarray_data_V_ce0       => FM_BBBB_L3PHID_enb,
      barrelFullMatches_15_dataarray_data_V_address0  => FM_BBBB_L3PHID_V_readaddr,
      barrelFullMatches_15_dataarray_data_V_q0        => FM_BBBB_L3PHID_V_dout,
      barrelFullMatches_15_nentries_0_V               => FM_BBBB_L3PHID_AV_dout_nent(0),
      barrelFullMatches_15_nentries_1_V               => FM_BBBB_L3PHID_AV_dout_nent(1),
      barrelFullMatches_16_dataarray_data_V_ce0       => FM_BBBB_L4PHIA_enb,
      barrelFullMatches_16_dataarray_data_V_address0  => FM_BBBB_L4PHIA_V_readaddr,
      barrelFullMatches_16_dataarray_data_V_q0        => FM_BBBB_L4PHIA_V_dout,
      barrelFullMatches_16_nentries_0_V               => FM_BBBB_L4PHIA_AV_dout_nent(0),
      barrelFullMatches_16_nentries_1_V               => FM_BBBB_L4PHIA_AV_dout_nent(1),
      barrelFullMatches_17_dataarray_data_V_ce0       => FM_BBBB_L4PHIB_enb,
      barrelFullMatches_17_dataarray_data_V_address0  => FM_BBBB_L4PHIB_V_readaddr,
      barrelFullMatches_17_dataarray_data_V_q0        => FM_BBBB_L4PHIB_V_dout,
      barrelFullMatches_17_nentries_0_V               => FM_BBBB_L4PHIB_AV_dout_nent(0),
      barrelFullMatches_17_nentries_1_V               => FM_BBBB_L4PHIB_AV_dout_nent(1),
      barrelFullMatches_18_dataarray_data_V_ce0       => FM_BBBB_L4PHIC_enb,
      barrelFullMatches_18_dataarray_data_V_address0  => FM_BBBB_L4PHIC_V_readaddr,
      barrelFullMatches_18_dataarray_data_V_q0        => FM_BBBB_L4PHIC_V_dout,
      barrelFullMatches_18_nentries_0_V               => FM_BBBB_L4PHIC_AV_dout_nent(0),
      barrelFullMatches_18_nentries_1_V               => FM_BBBB_L4PHIC_AV_dout_nent(1),
      barrelFullMatches_19_dataarray_data_V_ce0       => FM_BBBB_L4PHID_enb,
      barrelFullMatches_19_dataarray_data_V_address0  => FM_BBBB_L4PHID_V_readaddr,
      barrelFullMatches_19_dataarray_data_V_q0        => FM_BBBB_L4PHID_V_dout,
      barrelFullMatches_19_nentries_0_V               => FM_BBBB_L4PHID_AV_dout_nent(0),
      barrelFullMatches_19_nentries_1_V               => FM_BBBB_L4PHID_AV_dout_nent(1),
      barrelFullMatches_20_dataarray_data_V_ce0       => FM_BBBB_L5PHIA_enb,
      barrelFullMatches_20_dataarray_data_V_address0  => FM_BBBB_L5PHIA_V_readaddr,
      barrelFullMatches_20_dataarray_data_V_q0        => FM_BBBB_L5PHIA_V_dout,
      barrelFullMatches_20_nentries_0_V               => FM_BBBB_L5PHIA_AV_dout_nent(0),
      barrelFullMatches_20_nentries_1_V               => FM_BBBB_L5PHIA_AV_dout_nent(1),
      barrelFullMatches_21_dataarray_data_V_ce0       => FM_BBBB_L5PHIB_enb,
      barrelFullMatches_21_dataarray_data_V_address0  => FM_BBBB_L5PHIB_V_readaddr,
      barrelFullMatches_21_dataarray_data_V_q0        => FM_BBBB_L5PHIB_V_dout,
      barrelFullMatches_21_nentries_0_V               => FM_BBBB_L5PHIB_AV_dout_nent(0),
      barrelFullMatches_21_nentries_1_V               => FM_BBBB_L5PHIB_AV_dout_nent(1),
      barrelFullMatches_22_dataarray_data_V_ce0       => FM_BBBB_L5PHIC_enb,
      barrelFullMatches_22_dataarray_data_V_address0  => FM_BBBB_L5PHIC_V_readaddr,
      barrelFullMatches_22_dataarray_data_V_q0        => FM_BBBB_L5PHIC_V_dout,
      barrelFullMatches_22_nentries_0_V               => FM_BBBB_L5PHIC_AV_dout_nent(0),
      barrelFullMatches_22_nentries_1_V               => FM_BBBB_L5PHIC_AV_dout_nent(1),
      barrelFullMatches_23_dataarray_data_V_ce0       => FM_BBBB_L5PHID_enb,
      barrelFullMatches_23_dataarray_data_V_address0  => FM_BBBB_L5PHID_V_readaddr,
      barrelFullMatches_23_dataarray_data_V_q0        => FM_BBBB_L5PHID_V_dout,
      barrelFullMatches_23_nentries_0_V               => FM_BBBB_L5PHID_AV_dout_nent(0),
      barrelFullMatches_23_nentries_1_V               => FM_BBBB_L5PHID_AV_dout_nent(1),
      barrelFullMatches_24_dataarray_data_V_ce0       => FM_BBBB_L6PHIA_enb,
      barrelFullMatches_24_dataarray_data_V_address0  => FM_BBBB_L6PHIA_V_readaddr,
      barrelFullMatches_24_dataarray_data_V_q0        => FM_BBBB_L6PHIA_V_dout,
      barrelFullMatches_24_nentries_0_V               => FM_BBBB_L6PHIA_AV_dout_nent(0),
      barrelFullMatches_24_nentries_1_V               => FM_BBBB_L6PHIA_AV_dout_nent(1),
      barrelFullMatches_25_dataarray_data_V_ce0       => FM_BBBB_L6PHIB_enb,
      barrelFullMatches_25_dataarray_data_V_address0  => FM_BBBB_L6PHIB_V_readaddr,
      barrelFullMatches_25_dataarray_data_V_q0        => FM_BBBB_L6PHIB_V_dout,
      barrelFullMatches_25_nentries_0_V               => FM_BBBB_L6PHIB_AV_dout_nent(0),
      barrelFullMatches_25_nentries_1_V               => FM_BBBB_L6PHIB_AV_dout_nent(1),
      barrelFullMatches_26_dataarray_data_V_ce0       => FM_BBBB_L6PHIC_enb,
      barrelFullMatches_26_dataarray_data_V_address0  => FM_BBBB_L6PHIC_V_readaddr,
      barrelFullMatches_26_dataarray_data_V_q0        => FM_BBBB_L6PHIC_V_dout,
      barrelFullMatches_26_nentries_0_V               => FM_BBBB_L6PHIC_AV_dout_nent(0),
      barrelFullMatches_26_nentries_1_V               => FM_BBBB_L6PHIC_AV_dout_nent(1),
      barrelFullMatches_27_dataarray_data_V_ce0       => FM_BBBB_L6PHID_enb,
      barrelFullMatches_27_dataarray_data_V_address0  => FM_BBBB_L6PHID_V_readaddr,
      barrelFullMatches_27_dataarray_data_V_q0        => FM_BBBB_L6PHID_V_dout,
      barrelFullMatches_27_nentries_0_V               => FM_BBBB_L6PHID_AV_dout_nent(0),
      barrelFullMatches_27_nentries_1_V               => FM_BBBB_L6PHID_AV_dout_nent(1),
      diskFullMatches_0_dataarray_data_V_ce0       => FM_BBBB_D1PHIA_enb,
      diskFullMatches_0_dataarray_data_V_address0  => FM_BBBB_D1PHIA_V_readaddr,
      diskFullMatches_0_dataarray_data_V_q0        => FM_BBBB_D1PHIA_V_dout,
      diskFullMatches_0_nentries_0_V               => FM_BBBB_D1PHIA_AV_dout_nent(0),
      diskFullMatches_0_nentries_1_V               => FM_BBBB_D1PHIA_AV_dout_nent(1),
      diskFullMatches_1_dataarray_data_V_ce0       => FM_BBBB_D1PHIB_enb,
      diskFullMatches_1_dataarray_data_V_address0  => FM_BBBB_D1PHIB_V_readaddr,
      diskFullMatches_1_dataarray_data_V_q0        => FM_BBBB_D1PHIB_V_dout,
      diskFullMatches_1_nentries_0_V               => FM_BBBB_D1PHIB_AV_dout_nent(0),
      diskFullMatches_1_nentries_1_V               => FM_BBBB_D1PHIB_AV_dout_nent(1),
      diskFullMatches_2_dataarray_data_V_ce0       => FM_BBBB_D1PHIC_enb,
      diskFullMatches_2_dataarray_data_V_address0  => FM_BBBB_D1PHIC_V_readaddr,
      diskFullMatches_2_dataarray_data_V_q0        => FM_BBBB_D1PHIC_V_dout,
      diskFullMatches_2_nentries_0_V               => FM_BBBB_D1PHIC_AV_dout_nent(0),
      diskFullMatches_2_nentries_1_V               => FM_BBBB_D1PHIC_AV_dout_nent(1),
      diskFullMatches_3_dataarray_data_V_ce0       => FM_BBBB_D1PHID_enb,
      diskFullMatches_3_dataarray_data_V_address0  => FM_BBBB_D1PHID_V_readaddr,
      diskFullMatches_3_dataarray_data_V_q0        => FM_BBBB_D1PHID_V_dout,
      diskFullMatches_3_nentries_0_V               => FM_BBBB_D1PHID_AV_dout_nent(0),
      diskFullMatches_3_nentries_1_V               => FM_BBBB_D1PHID_AV_dout_nent(1),
      diskFullMatches_4_dataarray_data_V_ce0       => FM_BBBB_D2PHIA_enb,
      diskFullMatches_4_dataarray_data_V_address0  => FM_BBBB_D2PHIA_V_readaddr,
      diskFullMatches_4_dataarray_data_V_q0        => FM_BBBB_D2PHIA_V_dout,
      diskFullMatches_4_nentries_0_V               => FM_BBBB_D2PHIA_AV_dout_nent(0),
      diskFullMatches_4_nentries_1_V               => FM_BBBB_D2PHIA_AV_dout_nent(1),
      diskFullMatches_5_dataarray_data_V_ce0       => FM_BBBB_D2PHIB_enb,
      diskFullMatches_5_dataarray_data_V_address0  => FM_BBBB_D2PHIB_V_readaddr,
      diskFullMatches_5_dataarray_data_V_q0        => FM_BBBB_D2PHIB_V_dout,
      diskFullMatches_5_nentries_0_V               => FM_BBBB_D2PHIB_AV_dout_nent(0),
      diskFullMatches_5_nentries_1_V               => FM_BBBB_D2PHIB_AV_dout_nent(1),
      diskFullMatches_6_dataarray_data_V_ce0       => FM_BBBB_D2PHIC_enb,
      diskFullMatches_6_dataarray_data_V_address0  => FM_BBBB_D2PHIC_V_readaddr,
      diskFullMatches_6_dataarray_data_V_q0        => FM_BBBB_D2PHIC_V_dout,
      diskFullMatches_6_nentries_0_V               => FM_BBBB_D2PHIC_AV_dout_nent(0),
      diskFullMatches_6_nentries_1_V               => FM_BBBB_D2PHIC_AV_dout_nent(1),
      diskFullMatches_7_dataarray_data_V_ce0       => FM_BBBB_D2PHID_enb,
      diskFullMatches_7_dataarray_data_V_address0  => FM_BBBB_D2PHID_V_readaddr,
      diskFullMatches_7_dataarray_data_V_q0        => FM_BBBB_D2PHID_V_dout,
      diskFullMatches_7_nentries_0_V               => FM_BBBB_D2PHID_AV_dout_nent(0),
      diskFullMatches_7_nentries_1_V               => FM_BBBB_D2PHID_AV_dout_nent(1),
      diskFullMatches_8_dataarray_data_V_ce0       => FM_BBBB_D3PHIA_enb,
      diskFullMatches_8_dataarray_data_V_address0  => FM_BBBB_D3PHIA_V_readaddr,
      diskFullMatches_8_dataarray_data_V_q0        => FM_BBBB_D3PHIA_V_dout,
      diskFullMatches_8_nentries_0_V               => FM_BBBB_D3PHIA_AV_dout_nent(0),
      diskFullMatches_8_nentries_1_V               => FM_BBBB_D3PHIA_AV_dout_nent(1),
      diskFullMatches_9_dataarray_data_V_ce0       => FM_BBBB_D3PHIB_enb,
      diskFullMatches_9_dataarray_data_V_address0  => FM_BBBB_D3PHIB_V_readaddr,
      diskFullMatches_9_dataarray_data_V_q0        => FM_BBBB_D3PHIB_V_dout,
      diskFullMatches_9_nentries_0_V               => FM_BBBB_D3PHIB_AV_dout_nent(0),
      diskFullMatches_9_nentries_1_V               => FM_BBBB_D3PHIB_AV_dout_nent(1),
      diskFullMatches_10_dataarray_data_V_ce0       => FM_BBBB_D3PHIC_enb,
      diskFullMatches_10_dataarray_data_V_address0  => FM_BBBB_D3PHIC_V_readaddr,
      diskFullMatches_10_dataarray_data_V_q0        => FM_BBBB_D3PHIC_V_dout,
      diskFullMatches_10_nentries_0_V               => FM_BBBB_D3PHIC_AV_dout_nent(0),
      diskFullMatches_10_nentries_1_V               => FM_BBBB_D3PHIC_AV_dout_nent(1),
      diskFullMatches_11_dataarray_data_V_ce0       => FM_BBBB_D3PHID_enb,
      diskFullMatches_11_dataarray_data_V_address0  => FM_BBBB_D3PHID_V_readaddr,
      diskFullMatches_11_dataarray_data_V_q0        => FM_BBBB_D3PHID_V_dout,
      diskFullMatches_11_nentries_0_V               => FM_BBBB_D3PHID_AV_dout_nent(0),
      diskFullMatches_11_nentries_1_V               => FM_BBBB_D3PHID_AV_dout_nent(1),
      diskFullMatches_12_dataarray_data_V_ce0       => FM_BBBB_D4PHIA_enb,
      diskFullMatches_12_dataarray_data_V_address0  => FM_BBBB_D4PHIA_V_readaddr,
      diskFullMatches_12_dataarray_data_V_q0        => FM_BBBB_D4PHIA_V_dout,
      diskFullMatches_12_nentries_0_V               => FM_BBBB_D4PHIA_AV_dout_nent(0),
      diskFullMatches_12_nentries_1_V               => FM_BBBB_D4PHIA_AV_dout_nent(1),
      diskFullMatches_13_dataarray_data_V_ce0       => FM_BBBB_D4PHIB_enb,
      diskFullMatches_13_dataarray_data_V_address0  => FM_BBBB_D4PHIB_V_readaddr,
      diskFullMatches_13_dataarray_data_V_q0        => FM_BBBB_D4PHIB_V_dout,
      diskFullMatches_13_nentries_0_V               => FM_BBBB_D4PHIB_AV_dout_nent(0),
      diskFullMatches_13_nentries_1_V               => FM_BBBB_D4PHIB_AV_dout_nent(1),
      diskFullMatches_14_dataarray_data_V_ce0       => FM_BBBB_D4PHIC_enb,
      diskFullMatches_14_dataarray_data_V_address0  => FM_BBBB_D4PHIC_V_readaddr,
      diskFullMatches_14_dataarray_data_V_q0        => FM_BBBB_D4PHIC_V_dout,
      diskFullMatches_14_nentries_0_V               => FM_BBBB_D4PHIC_AV_dout_nent(0),
      diskFullMatches_14_nentries_1_V               => FM_BBBB_D4PHIC_AV_dout_nent(1),
      diskFullMatches_15_dataarray_data_V_ce0       => FM_BBBB_D4PHID_enb,
      diskFullMatches_15_dataarray_data_V_address0  => FM_BBBB_D4PHID_V_readaddr,
      diskFullMatches_15_dataarray_data_V_q0        => FM_BBBB_D4PHID_V_dout,
      diskFullMatches_15_nentries_0_V               => FM_BBBB_D4PHID_AV_dout_nent(0),
      diskFullMatches_15_nentries_1_V               => FM_BBBB_D4PHID_AV_dout_nent(1),
      diskFullMatches_16_dataarray_data_V_ce0       => FM_BBBB_D5PHIA_enb,
      diskFullMatches_16_dataarray_data_V_address0  => FM_BBBB_D5PHIA_V_readaddr,
      diskFullMatches_16_dataarray_data_V_q0        => FM_BBBB_D5PHIA_V_dout,
      diskFullMatches_16_nentries_0_V               => FM_BBBB_D5PHIA_AV_dout_nent(0),
      diskFullMatches_16_nentries_1_V               => FM_BBBB_D5PHIA_AV_dout_nent(1),
      diskFullMatches_17_dataarray_data_V_ce0       => FM_BBBB_D5PHIB_enb,
      diskFullMatches_17_dataarray_data_V_address0  => FM_BBBB_D5PHIB_V_readaddr,
      diskFullMatches_17_dataarray_data_V_q0        => FM_BBBB_D5PHIB_V_dout,
      diskFullMatches_17_nentries_0_V               => FM_BBBB_D5PHIB_AV_dout_nent(0),
      diskFullMatches_17_nentries_1_V               => FM_BBBB_D5PHIB_AV_dout_nent(1),
      diskFullMatches_18_dataarray_data_V_ce0       => FM_BBBB_D5PHIC_enb,
      diskFullMatches_18_dataarray_data_V_address0  => FM_BBBB_D5PHIC_V_readaddr,
      diskFullMatches_18_dataarray_data_V_q0        => FM_BBBB_D5PHIC_V_dout,
      diskFullMatches_18_nentries_0_V               => FM_BBBB_D5PHIC_AV_dout_nent(0),
      diskFullMatches_18_nentries_1_V               => FM_BBBB_D5PHIC_AV_dout_nent(1),
      diskFullMatches_19_dataarray_data_V_ce0       => FM_BBBB_D5PHID_enb,
      diskFullMatches_19_dataarray_data_V_address0  => FM_BBBB_D5PHID_V_readaddr,
      diskFullMatches_19_dataarray_data_V_q0        => FM_BBBB_D5PHID_V_dout,
      diskFullMatches_19_nentries_0_V               => FM_BBBB_D5PHID_AV_dout_nent(0),
      diskFullMatches_19_nentries_1_V               => FM_BBBB_D5PHID_AV_dout_nent(1),
      trackWord_V_din       => TW_BBBB_stream_AV_din,
      trackWord_V_full_n    => TW_BBBB_stream_A_full_neg,
      trackWord_V_write     => TW_BBBB_stream_A_write,
      barrelStubWords_0_V_din       => BW_BBBB_L1_stream_AV_din,
      barrelStubWords_0_V_full_n    => BW_BBBB_L1_stream_A_full_neg,
      barrelStubWords_0_V_write     => BW_BBBB_L1_stream_A_write,
      barrelStubWords_1_V_din       => BW_BBBB_L2_stream_AV_din,
      barrelStubWords_1_V_full_n    => BW_BBBB_L2_stream_A_full_neg,
      barrelStubWords_1_V_write     => BW_BBBB_L2_stream_A_write,
      barrelStubWords_2_V_din       => BW_BBBB_L3_stream_AV_din,
      barrelStubWords_2_V_full_n    => BW_BBBB_L3_stream_A_full_neg,
      barrelStubWords_2_V_write     => BW_BBBB_L3_stream_A_write,
      barrelStubWords_3_V_din       => BW_BBBB_L4_stream_AV_din,
      barrelStubWords_3_V_full_n    => BW_BBBB_L4_stream_A_full_neg,
      barrelStubWords_3_V_write     => BW_BBBB_L4_stream_A_write,
      barrelStubWords_4_V_din       => BW_BBBB_L5_stream_AV_din,
      barrelStubWords_4_V_full_n    => BW_BBBB_L5_stream_A_full_neg,
      barrelStubWords_4_V_write     => BW_BBBB_L5_stream_A_write,
      barrelStubWords_5_V_din       => BW_BBBB_L6_stream_AV_din,
      barrelStubWords_5_V_full_n    => BW_BBBB_L6_stream_A_full_neg,
      barrelStubWords_5_V_write     => BW_BBBB_L6_stream_A_write,
      diskStubWords_0_V_din       => DW_BBBB_D1_stream_AV_din,
      diskStubWords_0_V_full_n    => DW_BBBB_D1_stream_A_full_neg,
      diskStubWords_0_V_write     => DW_BBBB_D1_stream_A_write,
      diskStubWords_1_V_din       => DW_BBBB_D2_stream_AV_din,
      diskStubWords_1_V_full_n    => DW_BBBB_D2_stream_A_full_neg,
      diskStubWords_1_V_write     => DW_BBBB_D2_stream_A_write,
      diskStubWords_2_V_din       => DW_BBBB_D3_stream_AV_din,
      diskStubWords_2_V_full_n    => DW_BBBB_D3_stream_A_full_neg,
      diskStubWords_2_V_write     => DW_BBBB_D3_stream_A_write,
      diskStubWords_3_V_din       => DW_BBBB_D4_stream_AV_din,
      diskStubWords_3_V_full_n    => DW_BBBB_D4_stream_A_full_neg,
      diskStubWords_3_V_write     => DW_BBBB_D4_stream_A_write,
      diskStubWords_4_V_din       => DW_BBBB_D5_stream_AV_din,
      diskStubWords_4_V_full_n    => DW_BBBB_D5_stream_A_full_neg,
      diskStubWords_4_V_write     => DW_BBBB_D5_stream_A_write,
      done        => TB_BBBB_last_track,
      done_ap_vld => TB_BBBB_last_track_vld
  );

end rtl;
