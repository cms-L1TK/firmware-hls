--===========================================================================
--! @file
--! @brief Automatically generated top file for track finding.
--===========================================================================

--! Standard library
library ieee;
--! Standard package
use ieee.std_logic_1164.all;

--! User packages
use work.tf_pkg.all;


entity SectorProcessor is
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    en_proc    : in std_logic;
    bx_in_ProjectionRouter : in std_logic_vector(2 downto 0);
    bx_out_MatchCalculator : out std_logic_vector(2 downto 0);
    bx_out_MatchCalculator_vld : out std_logic;
    MatchCalculator_done   : out std_logic;
    TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L1L2XXG_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L1L2XXG_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXG_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L1L2XXG_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    VMSME_L3PHIC17n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC17n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC17n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC17n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC17n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC18n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC18n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC18n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC18n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC19n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC19n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC19n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC19n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC20n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC20n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC20n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC20n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC21n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC21n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC21n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC21n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC22n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC22n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC22n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC22n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC23n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC23n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC23n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC23n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_dataarray_data_V_wea       : in std_logic;
    VMSME_L3PHIC24n1_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    VMSME_L3PHIC24n1_dataarray_data_V_din       : in std_logic_vector(13 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_0_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_0_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_1_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_1_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_2_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_2_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_3_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_3_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_4_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_4_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_5_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_5_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_6_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_6_V_7_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_0_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_0_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_1_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_1_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_2_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_2_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_3_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_3_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_4_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_4_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_5_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_5_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_6_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_6_din  : in std_logic_vector(3 downto 0);
    VMSME_L3PHIC24n1_nentries_7_V_7_we   : in std_logic;
    VMSME_L3PHIC24n1_nentries_7_V_7_din  : in std_logic_vector(3 downto 0);
    TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L1L2XXH_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L1L2XXH_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXH_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L1L2XXH_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L1L2XXI_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L1L2XXI_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXI_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L1L2XXI_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L5L6XXC_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L5L6XXC_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXC_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L5L6XXC_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L5L6XXB_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L5L6XXB_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXB_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L5L6XXB_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L5L6XXD_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L5L6XXD_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L5L6XXD_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L5L6XXD_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_dataarray_data_V_wea       : in std_logic;
    AS_L3PHICn6_dataarray_data_V_writeaddr : in std_logic_vector(9 downto 0);
    AS_L3PHICn6_dataarray_data_V_din       : in std_logic_vector(35 downto 0);
    AS_L3PHICn6_nentries_0_V_we  : in std_logic;
    AS_L3PHICn6_nentries_0_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_1_V_we  : in std_logic;
    AS_L3PHICn6_nentries_1_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_2_V_we  : in std_logic;
    AS_L3PHICn6_nentries_2_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_3_V_we  : in std_logic;
    AS_L3PHICn6_nentries_3_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_4_V_we  : in std_logic;
    AS_L3PHICn6_nentries_4_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_5_V_we  : in std_logic;
    AS_L3PHICn6_nentries_5_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_6_V_we  : in std_logic;
    AS_L3PHICn6_nentries_6_V_din : in std_logic_vector(7 downto 0);
    AS_L3PHICn6_nentries_7_V_we  : in std_logic;
    AS_L3PHICn6_nentries_7_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_wea       : in std_logic;
    TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_writeaddr : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_din       : in std_logic_vector(59 downto 0);
    TPROJ_L1L2XXF_L3PHIC_nentries_0_V_we  : in std_logic;
    TPROJ_L1L2XXF_L3PHIC_nentries_0_V_din : in std_logic_vector(7 downto 0);
    TPROJ_L1L2XXF_L3PHIC_nentries_1_V_we  : in std_logic;
    TPROJ_L1L2XXF_L3PHIC_nentries_1_V_din : in std_logic_vector(7 downto 0);
    FM_L5L6_L3PHIC_dataarray_data_V_enb      : in std_logic;
    FM_L5L6_L3PHIC_dataarray_data_V_readaddr : in std_logic_vector(7 downto 0);
    FM_L5L6_L3PHIC_dataarray_data_V_dout     : out std_logic_vector(44 downto 0);
    FM_L5L6_L3PHIC_nentries_0_V_dout : out std_logic_vector(7 downto 0);
    FM_L5L6_L3PHIC_nentries_1_V_dout : out std_logic_vector(7 downto 0);
    FM_L1L2_L3PHIC_dataarray_data_V_enb      : in std_logic;
    FM_L1L2_L3PHIC_dataarray_data_V_readaddr : in std_logic_vector(7 downto 0);
    FM_L1L2_L3PHIC_dataarray_data_V_dout     : out std_logic_vector(44 downto 0);
    FM_L1L2_L3PHIC_nentries_0_V_dout : out std_logic_vector(7 downto 0);
    FM_L1L2_L3PHIC_nentries_1_V_dout : out std_logic_vector(7 downto 0)
);
end SectorProcessor;

architecture rtl of SectorProcessor is

  signal TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMSME_L3PHIC17n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC17n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC17n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC17n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC18n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC18n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC18n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC18n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC19n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC19n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC19n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC19n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC20n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC20n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC20n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC20n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC21n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC21n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC21n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC21n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC22n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC22n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC22n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC22n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC23n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC23n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC23n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC23n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);

  signal VMSME_L3PHIC24n1_dataarray_data_V_enb      : std_logic;
  signal VMSME_L3PHIC24n1_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal VMSME_L3PHIC24n1_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_0_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_1_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_2_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_3_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_4_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_5_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_6_V_7_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_0_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_1_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_2_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_3_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_4_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_5_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_6_dout : std_logic_vector(4 downto 0);
  signal VMSME_L3PHIC24n1_nentries_7_V_7_dout : std_logic_vector(4 downto 0);
  
  signal AS_L3PHICn6_dataarray_data_V_enb      : std_logic;
  signal AS_L3PHICn6_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal AS_L3PHICn6_dataarray_data_V_dout     : std_logic_vector(35 downto 0);
  signal AS_L3PHICn6_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_1_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_2_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_3_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_4_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_5_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_6_V_dout : std_logic_vector(7 downto 0);
  signal AS_L3PHICn6_nentries_7_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC17_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC17_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC17_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC17_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC17_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC17_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC17_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC17_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC17_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC17_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC17_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC17_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC18_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC18_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC18_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC18_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC18_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC18_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC18_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC18_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC18_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC18_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC18_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC18_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC19_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC19_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC19_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC19_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC19_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC19_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC19_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC19_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC19_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC19_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC19_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC19_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC20_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC20_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC20_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC20_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC20_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC20_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC20_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC20_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC20_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC20_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC20_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC20_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC21_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC21_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC21_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC21_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC21_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC21_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC21_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC21_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC21_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC21_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC21_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC21_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC22_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC22_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC22_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC22_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC22_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC22_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC22_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC22_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC22_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC22_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC22_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC22_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC23_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC23_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC23_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC23_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC23_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC23_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC23_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC23_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC23_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC23_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC23_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC23_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal VMPROJ_L3PHIC24_dataarray_data_V_wea       : std_logic;
  signal VMPROJ_L3PHIC24_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC24_dataarray_data_V_din       : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC24_nentries_0_V_we  : std_logic;
  signal VMPROJ_L3PHIC24_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC24_nentries_1_V_we  : std_logic;
  signal VMPROJ_L3PHIC24_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC24_dataarray_data_V_enb      : std_logic;
  signal VMPROJ_L3PHIC24_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC24_dataarray_data_V_dout     : std_logic_vector(20 downto 0);
  signal VMPROJ_L3PHIC24_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal VMPROJ_L3PHIC24_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC17_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC17_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC17_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC17_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC17_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC17_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC17_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC17_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC17_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC17_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC17_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC17_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC18_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC18_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC18_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC18_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC18_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC18_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC18_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC18_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC18_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC18_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC18_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC18_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC19_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC19_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC19_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC19_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC19_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC19_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC19_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC19_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC19_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC19_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC19_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC19_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC20_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC20_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC20_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC20_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC20_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC20_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC20_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC20_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC20_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC20_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC20_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC20_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC21_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC21_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC21_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC21_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC21_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC21_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC21_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC21_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC21_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC21_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC21_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC21_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC22_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC22_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC22_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC22_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC22_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC22_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC22_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC22_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC22_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC22_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC22_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC22_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC23_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC23_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC23_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC23_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC23_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC23_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC23_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC23_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC23_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC23_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC23_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC23_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal CM_L3PHIC24_dataarray_data_V_wea       : std_logic;
  signal CM_L3PHIC24_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC24_dataarray_data_V_din       : std_logic_vector(13 downto 0);
  signal CM_L3PHIC24_nentries_0_V_we  : std_logic;
  signal CM_L3PHIC24_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC24_nentries_1_V_we  : std_logic;
  signal CM_L3PHIC24_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal CM_L3PHIC24_dataarray_data_V_enb      : std_logic;
  signal CM_L3PHIC24_dataarray_data_V_readaddr : std_logic_vector(7 downto 0);
  signal CM_L3PHIC24_dataarray_data_V_dout     : std_logic_vector(13 downto 0);
  signal CM_L3PHIC24_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal CM_L3PHIC24_nentries_1_V_dout : std_logic_vector(7 downto 0);

  signal AP_L3PHIC_dataarray_data_V_wea       : std_logic;
  signal AP_L3PHIC_dataarray_data_V_writeaddr : std_logic_vector(9 downto 0);
  signal AP_L3PHIC_dataarray_data_V_din       : std_logic_vector(59 downto 0);
  signal AP_L3PHIC_nentries_0_V_we  : std_logic;
  signal AP_L3PHIC_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_1_V_we  : std_logic;
  signal AP_L3PHIC_nentries_1_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_2_V_we  : std_logic;
  signal AP_L3PHIC_nentries_2_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_3_V_we  : std_logic;
  signal AP_L3PHIC_nentries_3_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_4_V_we  : std_logic;
  signal AP_L3PHIC_nentries_4_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_5_V_we  : std_logic;
  signal AP_L3PHIC_nentries_5_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_6_V_we  : std_logic;
  signal AP_L3PHIC_nentries_6_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_7_V_we  : std_logic;
  signal AP_L3PHIC_nentries_7_V_din : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_dataarray_data_V_enb      : std_logic;
  signal AP_L3PHIC_dataarray_data_V_readaddr : std_logic_vector(9 downto 0);
  signal AP_L3PHIC_dataarray_data_V_dout     : std_logic_vector(59 downto 0);
  signal AP_L3PHIC_nentries_0_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_1_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_2_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_3_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_4_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_5_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_6_V_dout : std_logic_vector(7 downto 0);
  signal AP_L3PHIC_nentries_7_V_dout : std_logic_vector(7 downto 0);

  signal FM_L1L2_L3PHIC_dataarray_data_V_wea       : std_logic;
  signal FM_L1L2_L3PHIC_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal FM_L1L2_L3PHIC_dataarray_data_V_din       : std_logic_vector(44 downto 0);
  signal FM_L1L2_L3PHIC_nentries_0_V_we  : std_logic;
  signal FM_L1L2_L3PHIC_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal FM_L1L2_L3PHIC_nentries_1_V_we  : std_logic;
  signal FM_L1L2_L3PHIC_nentries_1_V_din : std_logic_vector(7 downto 0);

  signal FM_L5L6_L3PHIC_dataarray_data_V_wea       : std_logic;
  signal FM_L5L6_L3PHIC_dataarray_data_V_writeaddr : std_logic_vector(7 downto 0);
  signal FM_L5L6_L3PHIC_dataarray_data_V_din       : std_logic_vector(44 downto 0);
  signal FM_L5L6_L3PHIC_nentries_0_V_we  : std_logic;
  signal FM_L5L6_L3PHIC_nentries_0_V_din : std_logic_vector(7 downto 0);
  signal FM_L5L6_L3PHIC_nentries_1_V_we  : std_logic;
  signal FM_L5L6_L3PHIC_nentries_1_V_din : std_logic_vector(7 downto 0);

  signal ProjectionRouter_done : std_logic := '0';
  signal MatchEngine_start : std_logic := '0';
  signal bx_out_ProjectionRouter : std_logic_vector(2 downto 0);
  signal bx_out_ProjectionRouter_vld : std_logic;

  signal MatchEngine_done : std_logic := '0';
  signal MatchCalculator_start : std_logic := '0';
  signal bx_out_MatchEngine : std_logic_vector(2 downto 0);
  signal bx_out_MatchEngine_vld : std_logic;

begin

--  TPROJ_L1L2XXF_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L1L2XXF_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L1L2XXF_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L1L2XXF_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L1L2XXF_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L1L2XXG_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L1L2XXG_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L1L2XXG_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L1L2XXG_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L1L2XXG_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L1L2XXH_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L1L2XXH_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L1L2XXH_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L1L2XXH_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L1L2XXH_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L1L2XXI_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L1L2XXI_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L1L2XXI_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L1L2XXI_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L1L2XXI_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L1L2XXJ_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L5L6XXB_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L5L6XXB_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L5L6XXB_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L5L6XXB_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L5L6XXB_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L5L6XXC_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L5L6XXC_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L5L6XXC_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L5L6XXC_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L5L6XXC_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  TPROJ_L5L6XXD_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_wea,
--      addra     => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb,
--      addrb     => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => TPROJ_L5L6XXD_L3PHIC_nentries_0_V_we,
--      nent_i0  => TPROJ_L5L6XXD_L3PHIC_nentries_0_V_din,
--      nent_we1 => TPROJ_L5L6XXD_L3PHIC_nentries_1_V_we,
--      nent_i1  => TPROJ_L5L6XXD_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout,
--      nent_o1  => TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--VMSME_L3PHIC17n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC17n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC17n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC17n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC17n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC17n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC17n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC17n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC17n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC17n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC17n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC17n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC17n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC17n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC17n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC17n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC17n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC17n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC17n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC17n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC17n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC17n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC17n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC17n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC17n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC17n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC17n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC17n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC17n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC17n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC17n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC17n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC17n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC17n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC17n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC17n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC17n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC17n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC17n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC17n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC17n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC17n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC17n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC17n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC17n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC17n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC17n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC17n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC17n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC17n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC17n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC17n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC17n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC17n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC17n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC17n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC17n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC17n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC17n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC17n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC17n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC17n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC17n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC17n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC17n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC17n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC17n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC17n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC17n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC17n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC17n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC17n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC17n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC17n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC17n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC17n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC17n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC17n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC17n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC17n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC17n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC17n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC17n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC17n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC17n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC17n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC17n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC17n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC17n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC17n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC17n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC17n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC17n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC17n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC17n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC17n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC17n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC17n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC17n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC17n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC17n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC17n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC17n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC17n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC17n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC17n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC17n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC17n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC17n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC17n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC17n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC17n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC17n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC17n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC17n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC17n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC17n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC17n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC17n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC17n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC17n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC17n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC17n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC17n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC17n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC17n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC17n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC17n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC17n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC17n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC17n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC17n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC17n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC17n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC17n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC17n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC17n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC17n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC17n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC17n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC17n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC17n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC17n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC17n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC17n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC17n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC17n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC17n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC17n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC17n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC17n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC17n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC17n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC17n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC17n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC17n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC17n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC17n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC17n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC17n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC17n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC17n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC17n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC17n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC17n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC17n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC17n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC17n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC17n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC17n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC17n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC17n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC17n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC17n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC17n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC17n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC17n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC17n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC17n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC17n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC17n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC17n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC17n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC17n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC17n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC17n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC17n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC17n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC17n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC17n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC17n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC17n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC17n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC17n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC17n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC17n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC17n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC17n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC17n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC18n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC18n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC18n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC18n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC18n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC18n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC18n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC18n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC18n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC18n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC18n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC18n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC18n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC18n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC18n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC18n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC18n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC18n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC18n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC18n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC18n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC18n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC18n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC18n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC18n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC18n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC18n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC18n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC18n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC18n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC18n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC18n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC18n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC18n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC18n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC18n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC18n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC18n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC18n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC18n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC18n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC18n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC18n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC18n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC18n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC18n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC18n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC18n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC18n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC18n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC18n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC18n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC18n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC18n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC18n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC18n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC18n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC18n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC18n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC18n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC18n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC18n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC18n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC18n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC18n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC18n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC18n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC18n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC18n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC18n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC18n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC18n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC18n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC18n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC18n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC18n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC18n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC18n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC18n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC18n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC18n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC18n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC18n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC18n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC18n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC18n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC18n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC18n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC18n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC18n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC18n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC18n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC18n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC18n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC18n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC18n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC18n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC18n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC18n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC18n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC18n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC18n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC18n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC18n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC18n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC18n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC18n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC18n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC18n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC18n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC18n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC18n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC18n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC18n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC18n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC18n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC18n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC18n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC18n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC18n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC18n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC18n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC18n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC18n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC18n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC18n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC18n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC18n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC18n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC18n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC18n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC18n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC18n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC18n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC18n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC18n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC18n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC18n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC18n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC18n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC18n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC18n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC18n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC18n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC18n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC18n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC18n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC18n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC18n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC18n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC18n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC18n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC18n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC18n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC18n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC18n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC18n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC18n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC18n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC18n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC18n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC18n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC18n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC18n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC18n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC18n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC18n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC18n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC18n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC18n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC18n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC18n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC18n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC18n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC18n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC18n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC18n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC18n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC18n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC18n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC18n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC18n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC18n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC18n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC18n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC18n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC18n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC18n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC18n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC18n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC18n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC18n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC18n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC18n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC18n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC18n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC18n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC18n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC18n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC19n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC19n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC19n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC19n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC19n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC19n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC19n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC19n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC19n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC19n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC19n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC19n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC19n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC19n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC19n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC19n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC19n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC19n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC19n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC19n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC19n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC19n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC19n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC19n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC19n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC19n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC19n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC19n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC19n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC19n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC19n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC19n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC19n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC19n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC19n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC19n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC19n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC19n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC19n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC19n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC19n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC19n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC19n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC19n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC19n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC19n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC19n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC19n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC19n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC19n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC19n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC19n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC19n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC19n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC19n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC19n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC19n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC19n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC19n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC19n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC19n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC19n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC19n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC19n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC19n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC19n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC19n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC19n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC19n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC19n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC19n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC19n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC19n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC19n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC19n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC19n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC19n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC19n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC19n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC19n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC19n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC19n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC19n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC19n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC19n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC19n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC19n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC19n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC19n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC19n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC19n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC19n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC19n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC19n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC19n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC19n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC19n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC19n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC19n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC19n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC19n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC19n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC19n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC19n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC19n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC19n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC19n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC19n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC19n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC19n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC19n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC19n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC19n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC19n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC19n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC19n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC19n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC19n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC19n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC19n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC19n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC19n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC19n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC19n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC19n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC19n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC19n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC19n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC19n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC19n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC19n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC19n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC19n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC19n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC19n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC19n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC19n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC19n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC19n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC19n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC19n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC19n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC19n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC19n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC19n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC19n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC19n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC19n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC19n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC19n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC19n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC19n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC19n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC19n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC19n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC19n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC19n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC19n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC19n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC19n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC19n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC19n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC19n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC19n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC19n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC19n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC19n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC19n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC19n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC19n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC19n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC19n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC19n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC19n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC19n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC19n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC19n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC19n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC19n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC19n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC19n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC19n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC19n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC19n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC19n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC19n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC19n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC19n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC19n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC19n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC19n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC19n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC19n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC19n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC19n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC19n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC19n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC19n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC19n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC20n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC20n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC20n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC20n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC20n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC20n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC20n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC20n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC20n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC20n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC20n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC20n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC20n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC20n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC20n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC20n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC20n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC20n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC20n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC20n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC20n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC20n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC20n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC20n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC20n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC20n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC20n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC20n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC20n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC20n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC20n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC20n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC20n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC20n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC20n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC20n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC20n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC20n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC20n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC20n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC20n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC20n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC20n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC20n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC20n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC20n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC20n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC20n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC20n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC20n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC20n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC20n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC20n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC20n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC20n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC20n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC20n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC20n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC20n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC20n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC20n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC20n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC20n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC20n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC20n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC20n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC20n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC20n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC20n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC20n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC20n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC20n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC20n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC20n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC20n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC20n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC20n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC20n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC20n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC20n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC20n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC20n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC20n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC20n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC20n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC20n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC20n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC20n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC20n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC20n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC20n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC20n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC20n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC20n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC20n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC20n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC20n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC20n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC20n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC20n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC20n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC20n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC20n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC20n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC20n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC20n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC20n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC20n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC20n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC20n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC20n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC20n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC20n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC20n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC20n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC20n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC20n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC20n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC20n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC20n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC20n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC20n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC20n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC20n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC20n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC20n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC20n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC20n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC20n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC20n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC20n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC20n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC20n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC20n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC20n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC20n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC20n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC20n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC20n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC20n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC20n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC20n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC20n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC20n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC20n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC20n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC20n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC20n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC20n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC20n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC20n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC20n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC20n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC20n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC20n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC20n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC20n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC20n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC20n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC20n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC20n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC20n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC20n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC20n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC20n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC20n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC20n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC20n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC20n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC20n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC20n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC20n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC20n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC20n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC20n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC20n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC20n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC20n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC20n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC20n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC20n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC20n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC20n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC20n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC20n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC20n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC20n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC20n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC20n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC20n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC20n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC20n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC20n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC20n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC20n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC20n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC20n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC20n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC20n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC21n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC21n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC21n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC21n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC21n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC21n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC21n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC21n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC21n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC21n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC21n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC21n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC21n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC21n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC21n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC21n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC21n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC21n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC21n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC21n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC21n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC21n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC21n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC21n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC21n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC21n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC21n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC21n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC21n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC21n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC21n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC21n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC21n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC21n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC21n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC21n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC21n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC21n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC21n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC21n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC21n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC21n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC21n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC21n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC21n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC21n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC21n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC21n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC21n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC21n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC21n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC21n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC21n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC21n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC21n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC21n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC21n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC21n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC21n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC21n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC21n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC21n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC21n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC21n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC21n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC21n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC21n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC21n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC21n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC21n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC21n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC21n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC21n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC21n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC21n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC21n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC21n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC21n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC21n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC21n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC21n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC21n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC21n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC21n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC21n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC21n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC21n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC21n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC21n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC21n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC21n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC21n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC21n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC21n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC21n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC21n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC21n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC21n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC21n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC21n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC21n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC21n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC21n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC21n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC21n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC21n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC21n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC21n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC21n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC21n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC21n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC21n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC21n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC21n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC21n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC21n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC21n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC21n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC21n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC21n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC21n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC21n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC21n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC21n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC21n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC21n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC21n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC21n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC21n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC21n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC21n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC21n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC21n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC21n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC21n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC21n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC21n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC21n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC21n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC21n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC21n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC21n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC21n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC21n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC21n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC21n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC21n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC21n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC21n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC21n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC21n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC21n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC21n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC21n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC21n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC21n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC21n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC21n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC21n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC21n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC21n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC21n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC21n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC21n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC21n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC21n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC21n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC21n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC21n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC21n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC21n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC21n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC21n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC21n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC21n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC21n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC21n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC21n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC21n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC21n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC21n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC21n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC21n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC21n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC21n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC21n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC21n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC21n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC21n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC21n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC21n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC21n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC21n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC21n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC21n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC21n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC21n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC21n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC21n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC22n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC22n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC22n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC22n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC22n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC22n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC22n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC22n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC22n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC22n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC22n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC22n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC22n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC22n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC22n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC22n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC22n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC22n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC22n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC22n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC22n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC22n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC22n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC22n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC22n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC22n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC22n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC22n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC22n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC22n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC22n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC22n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC22n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC22n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC22n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC22n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC22n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC22n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC22n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC22n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC22n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC22n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC22n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC22n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC22n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC22n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC22n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC22n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC22n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC22n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC22n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC22n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC22n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC22n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC22n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC22n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC22n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC22n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC22n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC22n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC22n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC22n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC22n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC22n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC22n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC22n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC22n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC22n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC22n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC22n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC22n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC22n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC22n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC22n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC22n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC22n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC22n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC22n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC22n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC22n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC22n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC22n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC22n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC22n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC22n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC22n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC22n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC22n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC22n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC22n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC22n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC22n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC22n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC22n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC22n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC22n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC22n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC22n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC22n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC22n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC22n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC22n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC22n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC22n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC22n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC22n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC22n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC22n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC22n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC22n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC22n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC22n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC22n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC22n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC22n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC22n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC22n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC22n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC22n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC22n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC22n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC22n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC22n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC22n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC22n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC22n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC22n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC22n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC22n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC22n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC22n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC22n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC22n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC22n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC22n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC22n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC22n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC22n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC22n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC22n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC22n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC22n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC22n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC22n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC22n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC22n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC22n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC22n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC22n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC22n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC22n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC22n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC22n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC22n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC22n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC22n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC22n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC22n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC22n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC22n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC22n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC22n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC22n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC22n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC22n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC22n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC22n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC22n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC22n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC22n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC22n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC22n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC22n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC22n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC22n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC22n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC22n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC22n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC22n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC22n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC22n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC22n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC22n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC22n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC22n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC22n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC22n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC22n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC22n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC22n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC22n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC22n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC22n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC22n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC22n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC22n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC22n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC22n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC22n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC23n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC23n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC23n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC23n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC23n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC23n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC23n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC23n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC23n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC23n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC23n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC23n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC23n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC23n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC23n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC23n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC23n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC23n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC23n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC23n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC23n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC23n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC23n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC23n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC23n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC23n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC23n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC23n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC23n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC23n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC23n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC23n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC23n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC23n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC23n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC23n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC23n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC23n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC23n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC23n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC23n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC23n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC23n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC23n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC23n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC23n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC23n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC23n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC23n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC23n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC23n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC23n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC23n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC23n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC23n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC23n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC23n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC23n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC23n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC23n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC23n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC23n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC23n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC23n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC23n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC23n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC23n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC23n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC23n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC23n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC23n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC23n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC23n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC23n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC23n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC23n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC23n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC23n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC23n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC23n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC23n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC23n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC23n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC23n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC23n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC23n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC23n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC23n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC23n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC23n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC23n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC23n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC23n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC23n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC23n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC23n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC23n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC23n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC23n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC23n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC23n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC23n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC23n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC23n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC23n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC23n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC23n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC23n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC23n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC23n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC23n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC23n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC23n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC23n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC23n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC23n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC23n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC23n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC23n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC23n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC23n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC23n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC23n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC23n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC23n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC23n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC23n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC23n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC23n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC23n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC23n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC23n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC23n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC23n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC23n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC23n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC23n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC23n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC23n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC23n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC23n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC23n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC23n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC23n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC23n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC23n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC23n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC23n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC23n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC23n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC23n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC23n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC23n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC23n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC23n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC23n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC23n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC23n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC23n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC23n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC23n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC23n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC23n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC23n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC23n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC23n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC23n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC23n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC23n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC23n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC23n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC23n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC23n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC23n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC23n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC23n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC23n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC23n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC23n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC23n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC23n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC23n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC23n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC23n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC23n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC23n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC23n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC23n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC23n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC23n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC23n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC23n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC23n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC23n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC23n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC23n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC23n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC23n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC23n1_nentries_7_V_7_dout(3 downto 0)
--        );

--VMSME_L3PHIC24n1 : entity work.tf_mem_bin
--      generic map (
--        RAM_WIDTH       => 14,
--        RAM_DEPTH       => 1024,
--        INIT_FILE       => "",
--        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--        HEX             => 0       
--        )
--      port map (        
--        clka       => clk,
--        wea        => VMSME_L3PHIC24n1_dataarray_data_V_wea,
--        addra      => VMSME_L3PHIC24n1_dataarray_data_V_writeaddr(9 downto 0),
--        dina       => VMSME_L3PHIC24n1_dataarray_data_V_din,
--        nent_0_we0 =>  VMSME_L3PHIC24n1_nentries_0_V_0_we,
--        nent_0_i0  => VMSME_L3PHIC24n1_nentries_0_V_0_din,
--        nent_0_we1 =>  VMSME_L3PHIC24n1_nentries_0_V_1_we,
--        nent_0_i1  => VMSME_L3PHIC24n1_nentries_0_V_1_din,
--        nent_0_we2 =>  VMSME_L3PHIC24n1_nentries_0_V_2_we,
--        nent_0_i2  => VMSME_L3PHIC24n1_nentries_0_V_2_din,
--        nent_0_we3 =>  VMSME_L3PHIC24n1_nentries_0_V_3_we,
--        nent_0_i3  => VMSME_L3PHIC24n1_nentries_0_V_3_din,
--        nent_0_we4 =>  VMSME_L3PHIC24n1_nentries_0_V_4_we,
--        nent_0_i4  => VMSME_L3PHIC24n1_nentries_0_V_4_din,
--        nent_0_we5 =>  VMSME_L3PHIC24n1_nentries_0_V_5_we,
--        nent_0_i5  => VMSME_L3PHIC24n1_nentries_0_V_5_din,
--        nent_0_we6 =>  VMSME_L3PHIC24n1_nentries_0_V_6_we,
--        nent_0_i6  => VMSME_L3PHIC24n1_nentries_0_V_6_din,
--        nent_0_we7 =>  VMSME_L3PHIC24n1_nentries_0_V_7_we,
--        nent_0_i7  => VMSME_L3PHIC24n1_nentries_0_V_7_din,
--        nent_1_we0 =>  VMSME_L3PHIC24n1_nentries_1_V_0_we,
--        nent_1_i0  => VMSME_L3PHIC24n1_nentries_1_V_0_din,
--        nent_1_we1 =>  VMSME_L3PHIC24n1_nentries_1_V_1_we,
--        nent_1_i1  => VMSME_L3PHIC24n1_nentries_1_V_1_din,
--        nent_1_we2 =>  VMSME_L3PHIC24n1_nentries_1_V_2_we,
--        nent_1_i2  => VMSME_L3PHIC24n1_nentries_1_V_2_din,
--        nent_1_we3 =>  VMSME_L3PHIC24n1_nentries_1_V_3_we,
--        nent_1_i3  => VMSME_L3PHIC24n1_nentries_1_V_3_din,
--        nent_1_we4 =>  VMSME_L3PHIC24n1_nentries_1_V_4_we,
--        nent_1_i4  => VMSME_L3PHIC24n1_nentries_1_V_4_din,
--        nent_1_we5 =>  VMSME_L3PHIC24n1_nentries_1_V_5_we,
--        nent_1_i5  => VMSME_L3PHIC24n1_nentries_1_V_5_din,
--        nent_1_we6 =>  VMSME_L3PHIC24n1_nentries_1_V_6_we,
--        nent_1_i6  => VMSME_L3PHIC24n1_nentries_1_V_6_din,
--        nent_1_we7 =>  VMSME_L3PHIC24n1_nentries_1_V_7_we,
--        nent_1_i7  => VMSME_L3PHIC24n1_nentries_1_V_7_din,
--        nent_2_we0 =>  VMSME_L3PHIC24n1_nentries_2_V_0_we,
--        nent_2_i0  => VMSME_L3PHIC24n1_nentries_2_V_0_din,
--        nent_2_we1 =>  VMSME_L3PHIC24n1_nentries_2_V_1_we,
--        nent_2_i1  => VMSME_L3PHIC24n1_nentries_2_V_1_din,
--        nent_2_we2 =>  VMSME_L3PHIC24n1_nentries_2_V_2_we,
--        nent_2_i2  => VMSME_L3PHIC24n1_nentries_2_V_2_din,
--        nent_2_we3 =>  VMSME_L3PHIC24n1_nentries_2_V_3_we,
--        nent_2_i3  => VMSME_L3PHIC24n1_nentries_2_V_3_din,
--        nent_2_we4 =>  VMSME_L3PHIC24n1_nentries_2_V_4_we,
--        nent_2_i4  => VMSME_L3PHIC24n1_nentries_2_V_4_din,
--        nent_2_we5 =>  VMSME_L3PHIC24n1_nentries_2_V_5_we,
--        nent_2_i5  => VMSME_L3PHIC24n1_nentries_2_V_5_din,
--        nent_2_we6 =>  VMSME_L3PHIC24n1_nentries_2_V_6_we,
--        nent_2_i6  => VMSME_L3PHIC24n1_nentries_2_V_6_din,
--        nent_2_we7 =>  VMSME_L3PHIC24n1_nentries_2_V_7_we,
--        nent_2_i7  => VMSME_L3PHIC24n1_nentries_2_V_7_din,
--        nent_3_we0 =>  VMSME_L3PHIC24n1_nentries_3_V_0_we,
--        nent_3_i0  => VMSME_L3PHIC24n1_nentries_3_V_0_din,
--        nent_3_we1 =>  VMSME_L3PHIC24n1_nentries_3_V_1_we,
--        nent_3_i1  => VMSME_L3PHIC24n1_nentries_3_V_1_din,
--        nent_3_we2 =>  VMSME_L3PHIC24n1_nentries_3_V_2_we,
--        nent_3_i2  => VMSME_L3PHIC24n1_nentries_3_V_2_din,
--        nent_3_we3 =>  VMSME_L3PHIC24n1_nentries_3_V_3_we,
--        nent_3_i3  => VMSME_L3PHIC24n1_nentries_3_V_3_din,
--        nent_3_we4 =>  VMSME_L3PHIC24n1_nentries_3_V_4_we,
--        nent_3_i4  => VMSME_L3PHIC24n1_nentries_3_V_4_din,
--        nent_3_we5 =>  VMSME_L3PHIC24n1_nentries_3_V_5_we,
--        nent_3_i5  => VMSME_L3PHIC24n1_nentries_3_V_5_din,
--        nent_3_we6 =>  VMSME_L3PHIC24n1_nentries_3_V_6_we,
--        nent_3_i6  => VMSME_L3PHIC24n1_nentries_3_V_6_din,
--        nent_3_we7 =>  VMSME_L3PHIC24n1_nentries_3_V_7_we,
--        nent_3_i7  => VMSME_L3PHIC24n1_nentries_3_V_7_din,
--        nent_4_we0 =>  VMSME_L3PHIC24n1_nentries_4_V_0_we,
--        nent_4_i0  => VMSME_L3PHIC24n1_nentries_4_V_0_din,
--        nent_4_we1 =>  VMSME_L3PHIC24n1_nentries_4_V_1_we,
--        nent_4_i1  => VMSME_L3PHIC24n1_nentries_4_V_1_din,
--        nent_4_we2 =>  VMSME_L3PHIC24n1_nentries_4_V_2_we,
--        nent_4_i2  => VMSME_L3PHIC24n1_nentries_4_V_2_din,
--        nent_4_we3 =>  VMSME_L3PHIC24n1_nentries_4_V_3_we,
--        nent_4_i3  => VMSME_L3PHIC24n1_nentries_4_V_3_din,
--        nent_4_we4 =>  VMSME_L3PHIC24n1_nentries_4_V_4_we,
--        nent_4_i4  => VMSME_L3PHIC24n1_nentries_4_V_4_din,
--        nent_4_we5 =>  VMSME_L3PHIC24n1_nentries_4_V_5_we,
--        nent_4_i5  => VMSME_L3PHIC24n1_nentries_4_V_5_din,
--        nent_4_we6 =>  VMSME_L3PHIC24n1_nentries_4_V_6_we,
--        nent_4_i6  => VMSME_L3PHIC24n1_nentries_4_V_6_din,
--        nent_4_we7 =>  VMSME_L3PHIC24n1_nentries_4_V_7_we,
--        nent_4_i7  => VMSME_L3PHIC24n1_nentries_4_V_7_din,
--        nent_5_we0 =>  VMSME_L3PHIC24n1_nentries_5_V_0_we,
--        nent_5_i0  => VMSME_L3PHIC24n1_nentries_5_V_0_din,
--        nent_5_we1 =>  VMSME_L3PHIC24n1_nentries_5_V_1_we,
--        nent_5_i1  => VMSME_L3PHIC24n1_nentries_5_V_1_din,
--        nent_5_we2 =>  VMSME_L3PHIC24n1_nentries_5_V_2_we,
--        nent_5_i2  => VMSME_L3PHIC24n1_nentries_5_V_2_din,
--        nent_5_we3 =>  VMSME_L3PHIC24n1_nentries_5_V_3_we,
--        nent_5_i3  => VMSME_L3PHIC24n1_nentries_5_V_3_din,
--        nent_5_we4 =>  VMSME_L3PHIC24n1_nentries_5_V_4_we,
--        nent_5_i4  => VMSME_L3PHIC24n1_nentries_5_V_4_din,
--        nent_5_we5 =>  VMSME_L3PHIC24n1_nentries_5_V_5_we,
--        nent_5_i5  => VMSME_L3PHIC24n1_nentries_5_V_5_din,
--        nent_5_we6 =>  VMSME_L3PHIC24n1_nentries_5_V_6_we,
--        nent_5_i6  => VMSME_L3PHIC24n1_nentries_5_V_6_din,
--        nent_5_we7 =>  VMSME_L3PHIC24n1_nentries_5_V_7_we,
--        nent_5_i7  => VMSME_L3PHIC24n1_nentries_5_V_7_din,
--        nent_6_we0 =>  VMSME_L3PHIC24n1_nentries_6_V_0_we,
--        nent_6_i0  => VMSME_L3PHIC24n1_nentries_6_V_0_din,
--        nent_6_we1 =>  VMSME_L3PHIC24n1_nentries_6_V_1_we,
--        nent_6_i1  => VMSME_L3PHIC24n1_nentries_6_V_1_din,
--        nent_6_we2 =>  VMSME_L3PHIC24n1_nentries_6_V_2_we,
--        nent_6_i2  => VMSME_L3PHIC24n1_nentries_6_V_2_din,
--        nent_6_we3 =>  VMSME_L3PHIC24n1_nentries_6_V_3_we,
--        nent_6_i3  => VMSME_L3PHIC24n1_nentries_6_V_3_din,
--        nent_6_we4 =>  VMSME_L3PHIC24n1_nentries_6_V_4_we,
--        nent_6_i4  => VMSME_L3PHIC24n1_nentries_6_V_4_din,
--        nent_6_we5 =>  VMSME_L3PHIC24n1_nentries_6_V_5_we,
--        nent_6_i5  => VMSME_L3PHIC24n1_nentries_6_V_5_din,
--        nent_6_we6 =>  VMSME_L3PHIC24n1_nentries_6_V_6_we,
--        nent_6_i6  => VMSME_L3PHIC24n1_nentries_6_V_6_din,
--        nent_6_we7 =>  VMSME_L3PHIC24n1_nentries_6_V_7_we,
--        nent_6_i7  => VMSME_L3PHIC24n1_nentries_6_V_7_din,
--        nent_7_we0 =>  VMSME_L3PHIC24n1_nentries_7_V_0_we,
--        nent_7_i0  => VMSME_L3PHIC24n1_nentries_7_V_0_din,
--        nent_7_we1 =>  VMSME_L3PHIC24n1_nentries_7_V_1_we,
--        nent_7_i1  => VMSME_L3PHIC24n1_nentries_7_V_1_din,
--        nent_7_we2 =>  VMSME_L3PHIC24n1_nentries_7_V_2_we,
--        nent_7_i2  => VMSME_L3PHIC24n1_nentries_7_V_2_din,
--        nent_7_we3 =>  VMSME_L3PHIC24n1_nentries_7_V_3_we,
--        nent_7_i3  => VMSME_L3PHIC24n1_nentries_7_V_3_din,
--        nent_7_we4 =>  VMSME_L3PHIC24n1_nentries_7_V_4_we,
--        nent_7_i4  => VMSME_L3PHIC24n1_nentries_7_V_4_din,
--        nent_7_we5 =>  VMSME_L3PHIC24n1_nentries_7_V_5_we,
--        nent_7_i5  => VMSME_L3PHIC24n1_nentries_7_V_5_din,
--        nent_7_we6 =>  VMSME_L3PHIC24n1_nentries_7_V_6_we,
--        nent_7_i6  => VMSME_L3PHIC24n1_nentries_7_V_6_din,
--        nent_7_we7 =>  VMSME_L3PHIC24n1_nentries_7_V_7_we,
--        nent_7_i7  => VMSME_L3PHIC24n1_nentries_7_V_7_din,
--        clkb       => clk,
--        rstb       => '0',
--        regceb     => '1',
--        enb        => VMSME_L3PHIC24n1_dataarray_data_V_enb,
--        addrb      => VMSME_L3PHIC24n1_dataarray_data_V_readaddr,
--        doutb      => VMSME_L3PHIC24n1_dataarray_data_V_dout,
--        nent_0_o0  => VMSME_L3PHIC24n1_nentries_0_V_0_dout(3 downto 0),
--        nent_0_o1  => VMSME_L3PHIC24n1_nentries_0_V_1_dout(3 downto 0),
--        nent_0_o2  => VMSME_L3PHIC24n1_nentries_0_V_2_dout(3 downto 0),
--        nent_0_o3  => VMSME_L3PHIC24n1_nentries_0_V_3_dout(3 downto 0),
--        nent_0_o4  => VMSME_L3PHIC24n1_nentries_0_V_4_dout(3 downto 0),
--        nent_0_o5  => VMSME_L3PHIC24n1_nentries_0_V_5_dout(3 downto 0),
--        nent_0_o6  => VMSME_L3PHIC24n1_nentries_0_V_6_dout(3 downto 0),
--        nent_0_o7  => VMSME_L3PHIC24n1_nentries_0_V_7_dout(3 downto 0),
--        nent_1_o0  => VMSME_L3PHIC24n1_nentries_1_V_0_dout(3 downto 0),
--        nent_1_o1  => VMSME_L3PHIC24n1_nentries_1_V_1_dout(3 downto 0),
--        nent_1_o2  => VMSME_L3PHIC24n1_nentries_1_V_2_dout(3 downto 0),
--        nent_1_o3  => VMSME_L3PHIC24n1_nentries_1_V_3_dout(3 downto 0),
--        nent_1_o4  => VMSME_L3PHIC24n1_nentries_1_V_4_dout(3 downto 0),
--        nent_1_o5  => VMSME_L3PHIC24n1_nentries_1_V_5_dout(3 downto 0),
--        nent_1_o6  => VMSME_L3PHIC24n1_nentries_1_V_6_dout(3 downto 0),
--        nent_1_o7  => VMSME_L3PHIC24n1_nentries_1_V_7_dout(3 downto 0),
--        nent_2_o0  => VMSME_L3PHIC24n1_nentries_2_V_0_dout(3 downto 0),
--        nent_2_o1  => VMSME_L3PHIC24n1_nentries_2_V_1_dout(3 downto 0),
--        nent_2_o2  => VMSME_L3PHIC24n1_nentries_2_V_2_dout(3 downto 0),
--        nent_2_o3  => VMSME_L3PHIC24n1_nentries_2_V_3_dout(3 downto 0),
--        nent_2_o4  => VMSME_L3PHIC24n1_nentries_2_V_4_dout(3 downto 0),
--        nent_2_o5  => VMSME_L3PHIC24n1_nentries_2_V_5_dout(3 downto 0),
--        nent_2_o6  => VMSME_L3PHIC24n1_nentries_2_V_6_dout(3 downto 0),
--        nent_2_o7  => VMSME_L3PHIC24n1_nentries_2_V_7_dout(3 downto 0),
--        nent_3_o0  => VMSME_L3PHIC24n1_nentries_3_V_0_dout(3 downto 0),
--        nent_3_o1  => VMSME_L3PHIC24n1_nentries_3_V_1_dout(3 downto 0),
--        nent_3_o2  => VMSME_L3PHIC24n1_nentries_3_V_2_dout(3 downto 0),
--        nent_3_o3  => VMSME_L3PHIC24n1_nentries_3_V_3_dout(3 downto 0),
--        nent_3_o4  => VMSME_L3PHIC24n1_nentries_3_V_4_dout(3 downto 0),
--        nent_3_o5  => VMSME_L3PHIC24n1_nentries_3_V_5_dout(3 downto 0),
--        nent_3_o6  => VMSME_L3PHIC24n1_nentries_3_V_6_dout(3 downto 0),
--        nent_3_o7  => VMSME_L3PHIC24n1_nentries_3_V_7_dout(3 downto 0),
--        nent_4_o0  => VMSME_L3PHIC24n1_nentries_4_V_0_dout(3 downto 0),
--        nent_4_o1  => VMSME_L3PHIC24n1_nentries_4_V_1_dout(3 downto 0),
--        nent_4_o2  => VMSME_L3PHIC24n1_nentries_4_V_2_dout(3 downto 0),
--        nent_4_o3  => VMSME_L3PHIC24n1_nentries_4_V_3_dout(3 downto 0),
--        nent_4_o4  => VMSME_L3PHIC24n1_nentries_4_V_4_dout(3 downto 0),
--        nent_4_o5  => VMSME_L3PHIC24n1_nentries_4_V_5_dout(3 downto 0),
--        nent_4_o6  => VMSME_L3PHIC24n1_nentries_4_V_6_dout(3 downto 0),
--        nent_4_o7  => VMSME_L3PHIC24n1_nentries_4_V_7_dout(3 downto 0),
--        nent_5_o0  => VMSME_L3PHIC24n1_nentries_5_V_0_dout(3 downto 0),
--        nent_5_o1  => VMSME_L3PHIC24n1_nentries_5_V_1_dout(3 downto 0),
--        nent_5_o2  => VMSME_L3PHIC24n1_nentries_5_V_2_dout(3 downto 0),
--        nent_5_o3  => VMSME_L3PHIC24n1_nentries_5_V_3_dout(3 downto 0),
--        nent_5_o4  => VMSME_L3PHIC24n1_nentries_5_V_4_dout(3 downto 0),
--        nent_5_o5  => VMSME_L3PHIC24n1_nentries_5_V_5_dout(3 downto 0),
--        nent_5_o6  => VMSME_L3PHIC24n1_nentries_5_V_6_dout(3 downto 0),
--        nent_5_o7  => VMSME_L3PHIC24n1_nentries_5_V_7_dout(3 downto 0),
--        nent_6_o0  => VMSME_L3PHIC24n1_nentries_6_V_0_dout(3 downto 0),
--        nent_6_o1  => VMSME_L3PHIC24n1_nentries_6_V_1_dout(3 downto 0),
--        nent_6_o2  => VMSME_L3PHIC24n1_nentries_6_V_2_dout(3 downto 0),
--        nent_6_o3  => VMSME_L3PHIC24n1_nentries_6_V_3_dout(3 downto 0),
--        nent_6_o4  => VMSME_L3PHIC24n1_nentries_6_V_4_dout(3 downto 0),
--        nent_6_o5  => VMSME_L3PHIC24n1_nentries_6_V_5_dout(3 downto 0),
--        nent_6_o6  => VMSME_L3PHIC24n1_nentries_6_V_6_dout(3 downto 0),
--        nent_6_o7  => VMSME_L3PHIC24n1_nentries_6_V_7_dout(3 downto 0),
--        nent_7_o0  => VMSME_L3PHIC24n1_nentries_7_V_0_dout(3 downto 0),
--        nent_7_o1  => VMSME_L3PHIC24n1_nentries_7_V_1_dout(3 downto 0),
--        nent_7_o2  => VMSME_L3PHIC24n1_nentries_7_V_2_dout(3 downto 0),
--        nent_7_o3  => VMSME_L3PHIC24n1_nentries_7_V_3_dout(3 downto 0),
--        nent_7_o4  => VMSME_L3PHIC24n1_nentries_7_V_4_dout(3 downto 0),
--        nent_7_o5  => VMSME_L3PHIC24n1_nentries_7_V_5_dout(3 downto 0),
--        nent_7_o6  => VMSME_L3PHIC24n1_nentries_7_V_6_dout(3 downto 0),
--        nent_7_o7  => VMSME_L3PHIC24n1_nentries_7_V_7_dout(3 downto 0)
--        );


--  AS_L3PHICn6 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 36,
--      RAM_DEPTH       => 1024,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => AS_L3PHICn6_dataarray_data_V_wea,
--      addra     => AS_L3PHICn6_dataarray_data_V_writeaddr,
--      dina      => AS_L3PHICn6_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => AS_L3PHICn6_dataarray_data_V_enb,
--      addrb     => AS_L3PHICn6_dataarray_data_V_readaddr,
--      doutb     => AS_L3PHICn6_dataarray_data_V_dout,
--      nent_we0 => AS_L3PHICn6_nentries_0_V_we,
--      nent_i0  => AS_L3PHICn6_nentries_0_V_din,
--      nent_we1 => AS_L3PHICn6_nentries_1_V_we,
--      nent_i1  => AS_L3PHICn6_nentries_1_V_din,
--      nent_we2 => AS_L3PHICn6_nentries_2_V_we,
--      nent_i2  => AS_L3PHICn6_nentries_2_V_din,
--      nent_we3 => AS_L3PHICn6_nentries_3_V_we,
--      nent_i3  => AS_L3PHICn6_nentries_3_V_din,
--      nent_we4 => AS_L3PHICn6_nentries_4_V_we,
--      nent_i4  => AS_L3PHICn6_nentries_4_V_din,
--      nent_we5 => AS_L3PHICn6_nentries_5_V_we,
--      nent_i5  => AS_L3PHICn6_nentries_5_V_din,
--      nent_we6 => AS_L3PHICn6_nentries_6_V_we,
--      nent_i6  => AS_L3PHICn6_nentries_6_V_din,
--      nent_we7 => AS_L3PHICn6_nentries_7_V_we,
--      nent_i7  => AS_L3PHICn6_nentries_7_V_din,
--      nent_o0  => AS_L3PHICn6_nentries_0_V_dout,
--      nent_o1  => AS_L3PHICn6_nentries_1_V_dout,
--      nent_o2  => AS_L3PHICn6_nentries_2_V_dout,
--      nent_o3  => AS_L3PHICn6_nentries_3_V_dout,
--      nent_o4  => AS_L3PHICn6_nentries_4_V_dout,
--      nent_o5  => AS_L3PHICn6_nentries_5_V_dout,
--      nent_o6  => AS_L3PHICn6_nentries_6_V_dout,
--      nent_o7  => AS_L3PHICn6_nentries_7_V_dout
--  );


--  VMPROJ_L3PHIC17 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC17_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC17_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC17_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC17_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC17_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC17_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC17_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC17_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC17_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC17_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC17_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC17_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC18 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC18_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC18_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC18_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC18_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC18_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC18_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC18_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC18_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC18_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC18_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC18_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC18_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC19 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC19_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC19_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC19_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC19_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC19_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC19_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC19_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC19_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC19_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC19_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC19_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC19_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC20 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC20_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC20_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC20_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC20_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC20_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC20_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC20_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC20_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC20_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC20_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC20_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC20_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC21 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC21_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC21_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC21_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC21_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC21_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC21_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC21_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC21_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC21_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC21_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC21_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC21_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC22 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC22_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC22_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC22_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC22_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC22_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC22_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC22_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC22_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC22_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC22_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC22_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC22_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC23 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC23_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC23_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC23_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC23_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC23_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC23_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC23_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC23_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC23_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC23_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC23_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC23_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  VMPROJ_L3PHIC24 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 21,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => VMPROJ_L3PHIC24_dataarray_data_V_wea,
--      addra     => VMPROJ_L3PHIC24_dataarray_data_V_writeaddr,
--      dina      => VMPROJ_L3PHIC24_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => VMPROJ_L3PHIC24_dataarray_data_V_enb,
--      addrb     => VMPROJ_L3PHIC24_dataarray_data_V_readaddr,
--      doutb     => VMPROJ_L3PHIC24_dataarray_data_V_dout,
--      nent_we0 => VMPROJ_L3PHIC24_nentries_0_V_we,
--      nent_i0  => VMPROJ_L3PHIC24_nentries_0_V_din,
--      nent_we1 => VMPROJ_L3PHIC24_nentries_1_V_we,
--      nent_i1  => VMPROJ_L3PHIC24_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => VMPROJ_L3PHIC24_nentries_0_V_dout,
--      nent_o1  => VMPROJ_L3PHIC24_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC17 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC17_dataarray_data_V_wea,
--      addra     => CM_L3PHIC17_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC17_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC17_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC17_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC17_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC17_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC17_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC17_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC17_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC17_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC17_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC18 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC18_dataarray_data_V_wea,
--      addra     => CM_L3PHIC18_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC18_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC18_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC18_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC18_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC18_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC18_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC18_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC18_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC18_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC18_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC19 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC19_dataarray_data_V_wea,
--      addra     => CM_L3PHIC19_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC19_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC19_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC19_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC19_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC19_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC19_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC19_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC19_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC19_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC19_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC20 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC20_dataarray_data_V_wea,
--      addra     => CM_L3PHIC20_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC20_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC20_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC20_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC20_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC20_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC20_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC20_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC20_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC20_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC20_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC21 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC21_dataarray_data_V_wea,
--      addra     => CM_L3PHIC21_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC21_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC21_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC21_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC21_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC21_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC21_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC21_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC21_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC21_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC21_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC22 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC22_dataarray_data_V_wea,
--      addra     => CM_L3PHIC22_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC22_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC22_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC22_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC22_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC22_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC22_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC22_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC22_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC22_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC22_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC23 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC23_dataarray_data_V_wea,
--      addra     => CM_L3PHIC23_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC23_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC23_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC23_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC23_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC23_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC23_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC23_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC23_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC23_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC23_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  CM_L3PHIC24 : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 14,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => CM_L3PHIC24_dataarray_data_V_wea,
--      addra     => CM_L3PHIC24_dataarray_data_V_writeaddr,
--      dina      => CM_L3PHIC24_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => CM_L3PHIC24_dataarray_data_V_enb,
--      addrb     => CM_L3PHIC24_dataarray_data_V_readaddr,
--      doutb     => CM_L3PHIC24_dataarray_data_V_dout,
--      nent_we0 => CM_L3PHIC24_nentries_0_V_we,
--      nent_i0  => CM_L3PHIC24_nentries_0_V_din,
--      nent_we1 => CM_L3PHIC24_nentries_1_V_we,
--      nent_i1  => CM_L3PHIC24_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => CM_L3PHIC24_nentries_0_V_dout,
--      nent_o1  => CM_L3PHIC24_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  AP_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 60,
--      RAM_DEPTH       => 1024,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 1
--    )
--    port map (
--      clka      => clk,
--      wea       => AP_L3PHIC_dataarray_data_V_wea,
--      addra     => AP_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => AP_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => AP_L3PHIC_dataarray_data_V_enb,
--      addrb     => AP_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => AP_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => AP_L3PHIC_nentries_0_V_we,
--      nent_i0  => AP_L3PHIC_nentries_0_V_din,
--      nent_we1 => AP_L3PHIC_nentries_1_V_we,
--      nent_i1  => AP_L3PHIC_nentries_1_V_din,
--      nent_we2 => AP_L3PHIC_nentries_2_V_we,
--      nent_i2  => AP_L3PHIC_nentries_2_V_din,
--      nent_we3 => AP_L3PHIC_nentries_3_V_we,
--      nent_i3  => AP_L3PHIC_nentries_3_V_din,
--      nent_we4 => AP_L3PHIC_nentries_4_V_we,
--      nent_i4  => AP_L3PHIC_nentries_4_V_din,
--      nent_we5 => AP_L3PHIC_nentries_5_V_we,
--      nent_i5  => AP_L3PHIC_nentries_5_V_din,
--      nent_we6 => AP_L3PHIC_nentries_6_V_we,
--      nent_i6  => AP_L3PHIC_nentries_6_V_din,
--      nent_we7 => AP_L3PHIC_nentries_7_V_we,
--      nent_i7  => AP_L3PHIC_nentries_7_V_din,
--      nent_o0  => AP_L3PHIC_nentries_0_V_dout,
--      nent_o1  => AP_L3PHIC_nentries_1_V_dout,
--      nent_o2  => AP_L3PHIC_nentries_2_V_dout,
--      nent_o3  => AP_L3PHIC_nentries_3_V_dout,
--      nent_o4  => AP_L3PHIC_nentries_4_V_dout,
--      nent_o5  => AP_L3PHIC_nentries_5_V_dout,
--      nent_o6  => AP_L3PHIC_nentries_6_V_dout,
--      nent_o7  => AP_L3PHIC_nentries_7_V_dout
--  );


--  FM_L1L2_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 45,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => FM_L1L2_L3PHIC_dataarray_data_V_wea,
--      addra     => FM_L1L2_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => FM_L1L2_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => FM_L1L2_L3PHIC_dataarray_data_V_enb,
--      addrb     => FM_L1L2_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => FM_L1L2_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => FM_L1L2_L3PHIC_nentries_0_V_we,
--      nent_i0  => FM_L1L2_L3PHIC_nentries_0_V_din,
--      nent_we1 => FM_L1L2_L3PHIC_nentries_1_V_we,
--      nent_i1  => FM_L1L2_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => FM_L1L2_L3PHIC_nentries_0_V_dout,
--      nent_o1  => FM_L1L2_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );


--  FM_L5L6_L3PHIC : entity work.tf_mem
--    generic map (
--      RAM_WIDTH       => 45,
--      RAM_DEPTH       => 256,
--      INIT_FILE       => "",
--      RAM_PERFORMANCE => "HIGH_PERFORMANCE",
--      HEX             => 0
--    )
--    port map (
--      clka      => clk,
--      wea       => FM_L5L6_L3PHIC_dataarray_data_V_wea,
--      addra     => FM_L5L6_L3PHIC_dataarray_data_V_writeaddr,
--      dina      => FM_L5L6_L3PHIC_dataarray_data_V_din,
--      clkb      => clk,
--      rstb      => '0',
--      regceb    => '1',
--      enb       => FM_L5L6_L3PHIC_dataarray_data_V_enb,
--      addrb     => FM_L5L6_L3PHIC_dataarray_data_V_readaddr,
--      doutb     => FM_L5L6_L3PHIC_dataarray_data_V_dout,
--      nent_we0 => FM_L5L6_L3PHIC_nentries_0_V_we,
--      nent_i0  => FM_L5L6_L3PHIC_nentries_0_V_din,
--      nent_we1 => FM_L5L6_L3PHIC_nentries_1_V_we,
--      nent_i1  => FM_L5L6_L3PHIC_nentries_1_V_din,
--      nent_we2 => '0',
--      nent_i2  => (others=>'0'),
--      nent_we3 => '0',
--      nent_i3  => (others=>'0'),
--      nent_we4 => '0',
--      nent_i4  => (others=>'0'),
--      nent_we5 => '0',
--      nent_i5  => (others=>'0'),
--      nent_we6 => '0',
--      nent_i6  => (others=>'0'),
--      nent_we7 => '0',
--      nent_i7  => (others=>'0'),
--      nent_o0  => FM_L5L6_L3PHIC_nentries_0_V_dout,
--      nent_o1  => FM_L5L6_L3PHIC_nentries_1_V_dout,
--      nent_o2  => open,
--      nent_o3  => open,
--      nent_o4  => open,
--      nent_o5  => open,
--      nent_o6  => open,
--      nent_o7  => open
--  );

--  process(ProjectionRouter_done)
--  begin
--    if ProjectionRouter_done = '1' then MatchEngine_start <= '1'; end if;
--  end process;

--  PR_L3PHIC : entity work.PR_L3PHIC
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => en_proc,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => ProjectionRouter_done,
--      bx_V          => bx_in_ProjectionRouter,
--      bx_o_V        => bx_out_ProjectionRouter,
--      bx_o_V_ap_vld => bx_out_ProjectionRouter_vld,
--      projin_0_dataarray_data_V_ce0         => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb,
--      projin_0_dataarray_data_V_address0     => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr,
--      projin_0_dataarray_data_V_q0            => TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout,
--      projin_0_nentries_0_V        => TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_0_nentries_1_V        => TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_1_dataarray_data_V_ce0         => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb,
--      projin_1_dataarray_data_V_address0     => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr,
--      projin_1_dataarray_data_V_q0            => TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout,
--      projin_1_nentries_0_V        => TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_1_nentries_1_V        => TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_2_dataarray_data_V_ce0         => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb,
--      projin_2_dataarray_data_V_address0     => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr,
--      projin_2_dataarray_data_V_q0            => TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout,
--      projin_2_nentries_0_V        => TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_2_nentries_1_V        => TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_3_dataarray_data_V_ce0         => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb,
--      projin_3_dataarray_data_V_address0     => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr,
--      projin_3_dataarray_data_V_q0            => TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout,
--      projin_3_nentries_0_V        => TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_3_nentries_1_V        => TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_4_dataarray_data_V_ce0         => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb,
--      projin_4_dataarray_data_V_address0     => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr,
--      projin_4_dataarray_data_V_q0            => TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout,
--      projin_4_nentries_0_V        => TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_4_nentries_1_V        => TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_5_dataarray_data_V_ce0         => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb,
--      projin_5_dataarray_data_V_address0     => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr,
--      projin_5_dataarray_data_V_q0            => TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout,
--      projin_5_nentries_0_V        => TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_5_nentries_1_V        => TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_6_dataarray_data_V_ce0         => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb,
--      projin_6_dataarray_data_V_address0     => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr,
--      projin_6_dataarray_data_V_q0            => TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout,
--      projin_6_nentries_0_V        => TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_6_nentries_1_V        => TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout(6 downto 0),
--      projin_7_dataarray_data_V_ce0         => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb,
--      projin_7_dataarray_data_V_address0     => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr,
--      projin_7_dataarray_data_V_q0            => TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout,
--      projin_7_nentries_0_V        => TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout(6 downto 0),
--      projin_7_nentries_1_V        => TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout(6 downto 0),
--      allprojout_dataarray_data_V_ce0         => open,
--      allprojout_dataarray_data_V_we0         => AP_L3PHIC_dataarray_data_V_wea,
--      allprojout_dataarray_data_V_address0    => AP_L3PHIC_dataarray_data_V_writeaddr,
--      allprojout_dataarray_data_V_d0          => AP_L3PHIC_dataarray_data_V_din,
--      vmprojout_0_dataarray_data_V_ce0         => open,
--      vmprojout_0_dataarray_data_V_we0         => VMPROJ_L3PHIC17_dataarray_data_V_wea,
--      vmprojout_0_dataarray_data_V_address0    => VMPROJ_L3PHIC17_dataarray_data_V_writeaddr,
--      vmprojout_0_dataarray_data_V_d0          => VMPROJ_L3PHIC17_dataarray_data_V_din,
--      vmprojout_1_dataarray_data_V_ce0         => open,
--      vmprojout_1_dataarray_data_V_we0         => VMPROJ_L3PHIC18_dataarray_data_V_wea,
--      vmprojout_1_dataarray_data_V_address0    => VMPROJ_L3PHIC18_dataarray_data_V_writeaddr,
--      vmprojout_1_dataarray_data_V_d0          => VMPROJ_L3PHIC18_dataarray_data_V_din,
--      vmprojout_2_dataarray_data_V_ce0         => open,
--      vmprojout_2_dataarray_data_V_we0         => VMPROJ_L3PHIC19_dataarray_data_V_wea,
--      vmprojout_2_dataarray_data_V_address0    => VMPROJ_L3PHIC19_dataarray_data_V_writeaddr,
--      vmprojout_2_dataarray_data_V_d0          => VMPROJ_L3PHIC19_dataarray_data_V_din,
--      vmprojout_3_dataarray_data_V_ce0         => open,
--      vmprojout_3_dataarray_data_V_we0         => VMPROJ_L3PHIC20_dataarray_data_V_wea,
--      vmprojout_3_dataarray_data_V_address0    => VMPROJ_L3PHIC20_dataarray_data_V_writeaddr,
--      vmprojout_3_dataarray_data_V_d0          => VMPROJ_L3PHIC20_dataarray_data_V_din,
--      vmprojout_4_dataarray_data_V_ce0         => open,
--      vmprojout_4_dataarray_data_V_we0         => VMPROJ_L3PHIC21_dataarray_data_V_wea,
--      vmprojout_4_dataarray_data_V_address0    => VMPROJ_L3PHIC21_dataarray_data_V_writeaddr,
--      vmprojout_4_dataarray_data_V_d0          => VMPROJ_L3PHIC21_dataarray_data_V_din,
--      vmprojout_5_dataarray_data_V_ce0         => open,
--      vmprojout_5_dataarray_data_V_we0         => VMPROJ_L3PHIC22_dataarray_data_V_wea,
--      vmprojout_5_dataarray_data_V_address0    => VMPROJ_L3PHIC22_dataarray_data_V_writeaddr,
--      vmprojout_5_dataarray_data_V_d0          => VMPROJ_L3PHIC22_dataarray_data_V_din,
--      vmprojout_6_dataarray_data_V_ce0         => open,
--      vmprojout_6_dataarray_data_V_we0         => VMPROJ_L3PHIC23_dataarray_data_V_wea,
--      vmprojout_6_dataarray_data_V_address0    => VMPROJ_L3PHIC23_dataarray_data_V_writeaddr,
--      vmprojout_6_dataarray_data_V_d0          => VMPROJ_L3PHIC23_dataarray_data_V_din,
--      vmprojout_7_dataarray_data_V_ce0         => open,
--      vmprojout_7_dataarray_data_V_we0         => VMPROJ_L3PHIC24_dataarray_data_V_wea,
--      vmprojout_7_dataarray_data_V_address0    => VMPROJ_L3PHIC24_dataarray_data_V_writeaddr,
--      vmprojout_7_dataarray_data_V_d0          => VMPROJ_L3PHIC24_dataarray_data_V_din  );

--  process(MatchEngine_done)
--  begin
--    if MatchEngine_done = '1' then MatchCalculator_start <= '1'; end if;
--  end process;

--  ME_L3PHIC17 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC17n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC17n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC17n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC17n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC17n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC17n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC17n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC17n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC17n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC17n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC17n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC17n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC17n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC17n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC17n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC17n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC17n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC17n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC17n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC17n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC17n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC17n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC17n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC17n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC17n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC17n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC17n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC17n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC17n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC17n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC17n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC17n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC17n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC17n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC17n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC17n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC17n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC17n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC17n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC17n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC17n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC17n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC17n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC17n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC17n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC17n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC17n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC17n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC17n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC17n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC17n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC17n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC17n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC17n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC17n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC17n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC17n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC17n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC17n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC17n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC17n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC17n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC17n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC17n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC17n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC17n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC17n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC17_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC17_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC17_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC17_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC17_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC17_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC17_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC17_dataarray_data_V_din  );

--  ME_L3PHIC18 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC18n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC18n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC18n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC18n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC18n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC18n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC18n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC18n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC18n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC18n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC18n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC18n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC18n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC18n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC18n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC18n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC18n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC18n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC18n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC18n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC18n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC18n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC18n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC18n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC18n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC18n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC18n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC18n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC18n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC18n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC18n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC18n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC18n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC18n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC18n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC18n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC18n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC18n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC18n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC18n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC18n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC18n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC18n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC18n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC18n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC18n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC18n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC18n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC18n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC18n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC18n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC18n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC18n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC18n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC18n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC18n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC18n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC18n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC18n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC18n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC18n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC18n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC18n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC18n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC18n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC18n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC18n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC18_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC18_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC18_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC18_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC18_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC18_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC18_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC18_dataarray_data_V_din  );

--  ME_L3PHIC19 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC19n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC19n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC19n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC19n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC19n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC19n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC19n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC19n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC19n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC19n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC19n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC19n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC19n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC19n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC19n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC19n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC19n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC19n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC19n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC19n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC19n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC19n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC19n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC19n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC19n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC19n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC19n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC19n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC19n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC19n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC19n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC19n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC19n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC19n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC19n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC19n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC19n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC19n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC19n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC19n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC19n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC19n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC19n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC19n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC19n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC19n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC19n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC19n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC19n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC19n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC19n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC19n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC19n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC19n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC19n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC19n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC19n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC19n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC19n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC19n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC19n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC19n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC19n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC19n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC19n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC19n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC19n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC19_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC19_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC19_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC19_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC19_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC19_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC19_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC19_dataarray_data_V_din  );

--  ME_L3PHIC20 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC20n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC20n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC20n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC20n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC20n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC20n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC20n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC20n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC20n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC20n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC20n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC20n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC20n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC20n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC20n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC20n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC20n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC20n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC20n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC20n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC20n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC20n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC20n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC20n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC20n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC20n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC20n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC20n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC20n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC20n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC20n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC20n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC20n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC20n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC20n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC20n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC20n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC20n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC20n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC20n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC20n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC20n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC20n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC20n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC20n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC20n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC20n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC20n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC20n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC20n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC20n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC20n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC20n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC20n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC20n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC20n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC20n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC20n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC20n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC20n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC20n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC20n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC20n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC20n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC20n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC20n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC20n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC20_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC20_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC20_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC20_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC20_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC20_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC20_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC20_dataarray_data_V_din  );

--  ME_L3PHIC21 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC21n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC21n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC21n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC21n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC21n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC21n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC21n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC21n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC21n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC21n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC21n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC21n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC21n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC21n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC21n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC21n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC21n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC21n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC21n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC21n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC21n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC21n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC21n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC21n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC21n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC21n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC21n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC21n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC21n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC21n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC21n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC21n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC21n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC21n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC21n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC21n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC21n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC21n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC21n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC21n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC21n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC21n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC21n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC21n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC21n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC21n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC21n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC21n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC21n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC21n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC21n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC21n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC21n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC21n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC21n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC21n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC21n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC21n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC21n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC21n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC21n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC21n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC21n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC21n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC21n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC21n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC21n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC21_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC21_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC21_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC21_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC21_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC21_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC21_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC21_dataarray_data_V_din  );

--  ME_L3PHIC22 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC22n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC22n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC22n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC22n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC22n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC22n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC22n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC22n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC22n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC22n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC22n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC22n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC22n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC22n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC22n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC22n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC22n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC22n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC22n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC22n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC22n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC22n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC22n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC22n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC22n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC22n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC22n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC22n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC22n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC22n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC22n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC22n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC22n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC22n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC22n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC22n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC22n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC22n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC22n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC22n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC22n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC22n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC22n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC22n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC22n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC22n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC22n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC22n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC22n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC22n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC22n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC22n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC22n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC22n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC22n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC22n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC22n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC22n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC22n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC22n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC22n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC22n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC22n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC22n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC22n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC22n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC22n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC22_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC22_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC22_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC22_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC22_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC22_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC22_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC22_dataarray_data_V_din  );

--  ME_L3PHIC23 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC23n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC23n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC23n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC23n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC23n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC23n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC23n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC23n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC23n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC23n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC23n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC23n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC23n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC23n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC23n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC23n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC23n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC23n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC23n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC23n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC23n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC23n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC23n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC23n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC23n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC23n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC23n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC23n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC23n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC23n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC23n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC23n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC23n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC23n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC23n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC23n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC23n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC23n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC23n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC23n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC23n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC23n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC23n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC23n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC23n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC23n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC23n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC23n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC23n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC23n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC23n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC23n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC23n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC23n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC23n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC23n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC23n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC23n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC23n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC23n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC23n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC23n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC23n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC23n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC23n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC23n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC23n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC23_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC23_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC23_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC23_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC23_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC23_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC23_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC23_dataarray_data_V_din  );

--  ME_L3PHIC24 : entity work.MatchEngineTopL3_0 
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchEngine_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchEngine_done,
--      bx_V          => bx_out_ProjectionRouter,
--      bx_o_V        => bx_out_MatchEngine,
--      bx_o_V_ap_vld => bx_out_MatchEngine_vld,
--      inputStubData_dataarray_data_V_ce0         => VMSME_L3PHIC24n1_dataarray_data_V_enb,
--      inputStubData_dataarray_data_V_address0     => VMSME_L3PHIC24n1_dataarray_data_V_readaddr,
--      inputStubData_dataarray_data_V_q0            => VMSME_L3PHIC24n1_dataarray_data_V_dout(12 downto 0),
--      inputStubData_nentries_0_V_0 => VMSME_L3PHIC24n1_nentries_0_V_0_dout,
--      inputStubData_nentries_0_V_1 => VMSME_L3PHIC24n1_nentries_0_V_1_dout,
--      inputStubData_nentries_0_V_2 => VMSME_L3PHIC24n1_nentries_0_V_2_dout,
--      inputStubData_nentries_0_V_3 => VMSME_L3PHIC24n1_nentries_0_V_3_dout,
--      inputStubData_nentries_0_V_4 => VMSME_L3PHIC24n1_nentries_0_V_4_dout,
--      inputStubData_nentries_0_V_5 => VMSME_L3PHIC24n1_nentries_0_V_5_dout,
--      inputStubData_nentries_0_V_6 => VMSME_L3PHIC24n1_nentries_0_V_6_dout,
--      inputStubData_nentries_0_V_7 => VMSME_L3PHIC24n1_nentries_0_V_7_dout,
--      inputStubData_nentries_1_V_0 => VMSME_L3PHIC24n1_nentries_1_V_0_dout,
--      inputStubData_nentries_1_V_1 => VMSME_L3PHIC24n1_nentries_1_V_1_dout,
--      inputStubData_nentries_1_V_2 => VMSME_L3PHIC24n1_nentries_1_V_2_dout,
--      inputStubData_nentries_1_V_3 => VMSME_L3PHIC24n1_nentries_1_V_3_dout,
--      inputStubData_nentries_1_V_4 => VMSME_L3PHIC24n1_nentries_1_V_4_dout,
--      inputStubData_nentries_1_V_5 => VMSME_L3PHIC24n1_nentries_1_V_5_dout,
--      inputStubData_nentries_1_V_6 => VMSME_L3PHIC24n1_nentries_1_V_6_dout,
--      inputStubData_nentries_1_V_7 => VMSME_L3PHIC24n1_nentries_1_V_7_dout,
--      inputStubData_nentries_2_V_0 => VMSME_L3PHIC24n1_nentries_2_V_0_dout,
--      inputStubData_nentries_2_V_1 => VMSME_L3PHIC24n1_nentries_2_V_1_dout,
--      inputStubData_nentries_2_V_2 => VMSME_L3PHIC24n1_nentries_2_V_2_dout,
--      inputStubData_nentries_2_V_3 => VMSME_L3PHIC24n1_nentries_2_V_3_dout,
--      inputStubData_nentries_2_V_4 => VMSME_L3PHIC24n1_nentries_2_V_4_dout,
--      inputStubData_nentries_2_V_5 => VMSME_L3PHIC24n1_nentries_2_V_5_dout,
--      inputStubData_nentries_2_V_6 => VMSME_L3PHIC24n1_nentries_2_V_6_dout,
--      inputStubData_nentries_2_V_7 => VMSME_L3PHIC24n1_nentries_2_V_7_dout,
--      inputStubData_nentries_3_V_0 => VMSME_L3PHIC24n1_nentries_3_V_0_dout,
--      inputStubData_nentries_3_V_1 => VMSME_L3PHIC24n1_nentries_3_V_1_dout,
--      inputStubData_nentries_3_V_2 => VMSME_L3PHIC24n1_nentries_3_V_2_dout,
--      inputStubData_nentries_3_V_3 => VMSME_L3PHIC24n1_nentries_3_V_3_dout,
--      inputStubData_nentries_3_V_4 => VMSME_L3PHIC24n1_nentries_3_V_4_dout,
--      inputStubData_nentries_3_V_5 => VMSME_L3PHIC24n1_nentries_3_V_5_dout,
--      inputStubData_nentries_3_V_6 => VMSME_L3PHIC24n1_nentries_3_V_6_dout,
--      inputStubData_nentries_3_V_7 => VMSME_L3PHIC24n1_nentries_3_V_7_dout,
--      inputStubData_nentries_4_V_0 => VMSME_L3PHIC24n1_nentries_4_V_0_dout,
--      inputStubData_nentries_4_V_1 => VMSME_L3PHIC24n1_nentries_4_V_1_dout,
--      inputStubData_nentries_4_V_2 => VMSME_L3PHIC24n1_nentries_4_V_2_dout,
--      inputStubData_nentries_4_V_3 => VMSME_L3PHIC24n1_nentries_4_V_3_dout,
--      inputStubData_nentries_4_V_4 => VMSME_L3PHIC24n1_nentries_4_V_4_dout,
--      inputStubData_nentries_4_V_5 => VMSME_L3PHIC24n1_nentries_4_V_5_dout,
--      inputStubData_nentries_4_V_6 => VMSME_L3PHIC24n1_nentries_4_V_6_dout,
--      inputStubData_nentries_4_V_7 => VMSME_L3PHIC24n1_nentries_4_V_7_dout,
--      inputStubData_nentries_5_V_0 => VMSME_L3PHIC24n1_nentries_5_V_0_dout,
--      inputStubData_nentries_5_V_1 => VMSME_L3PHIC24n1_nentries_5_V_1_dout,
--      inputStubData_nentries_5_V_2 => VMSME_L3PHIC24n1_nentries_5_V_2_dout,
--      inputStubData_nentries_5_V_3 => VMSME_L3PHIC24n1_nentries_5_V_3_dout,
--      inputStubData_nentries_5_V_4 => VMSME_L3PHIC24n1_nentries_5_V_4_dout,
--      inputStubData_nentries_5_V_5 => VMSME_L3PHIC24n1_nentries_5_V_5_dout,
--      inputStubData_nentries_5_V_6 => VMSME_L3PHIC24n1_nentries_5_V_6_dout,
--      inputStubData_nentries_5_V_7 => VMSME_L3PHIC24n1_nentries_5_V_7_dout,
--      inputStubData_nentries_6_V_0 => VMSME_L3PHIC24n1_nentries_6_V_0_dout,
--      inputStubData_nentries_6_V_1 => VMSME_L3PHIC24n1_nentries_6_V_1_dout,
--      inputStubData_nentries_6_V_2 => VMSME_L3PHIC24n1_nentries_6_V_2_dout,
--      inputStubData_nentries_6_V_3 => VMSME_L3PHIC24n1_nentries_6_V_3_dout,
--      inputStubData_nentries_6_V_4 => VMSME_L3PHIC24n1_nentries_6_V_4_dout,
--      inputStubData_nentries_6_V_5 => VMSME_L3PHIC24n1_nentries_6_V_5_dout,
--      inputStubData_nentries_6_V_6 => VMSME_L3PHIC24n1_nentries_6_V_6_dout,
--      inputStubData_nentries_6_V_7 => VMSME_L3PHIC24n1_nentries_6_V_7_dout,
--      inputStubData_nentries_7_V_0 => VMSME_L3PHIC24n1_nentries_7_V_0_dout,
--      inputStubData_nentries_7_V_1 => VMSME_L3PHIC24n1_nentries_7_V_1_dout,
--      inputStubData_nentries_7_V_2 => VMSME_L3PHIC24n1_nentries_7_V_2_dout,
--      inputStubData_nentries_7_V_3 => VMSME_L3PHIC24n1_nentries_7_V_3_dout,
--      inputStubData_nentries_7_V_4 => VMSME_L3PHIC24n1_nentries_7_V_4_dout,
--      inputStubData_nentries_7_V_5 => VMSME_L3PHIC24n1_nentries_7_V_5_dout,
--      inputStubData_nentries_7_V_6 => VMSME_L3PHIC24n1_nentries_7_V_6_dout,
--      inputStubData_nentries_7_V_7 => VMSME_L3PHIC24n1_nentries_7_V_7_dout,
--      inputProjectionData_dataarray_data_V_ce0         => VMPROJ_L3PHIC24_dataarray_data_V_enb,
--      inputProjectionData_dataarray_data_V_address0     => VMPROJ_L3PHIC24_dataarray_data_V_readaddr,
--      inputProjectionData_dataarray_data_V_q0            => VMPROJ_L3PHIC24_dataarray_data_V_dout,
--      inputProjectionData_nentries_0_V        => VMPROJ_L3PHIC24_nentries_0_V_dout(6 downto 0),
--      inputProjectionData_nentries_1_V        => VMPROJ_L3PHIC24_nentries_1_V_dout(6 downto 0),
--      outputCandidateMatch_dataarray_data_V_ce0         => open,
--      outputCandidateMatch_dataarray_data_V_we0         => CM_L3PHIC24_dataarray_data_V_wea,
--      outputCandidateMatch_dataarray_data_V_address0    => CM_L3PHIC24_dataarray_data_V_writeaddr,
--      outputCandidateMatch_dataarray_data_V_d0          => CM_L3PHIC24_dataarray_data_V_din  );

--  MC_L3PHIC : entity work.MC_L3PHIC
--    port map (
--      ap_clk   => clk,
--      ap_rst   => reset,
--      ap_start => MatchCalculator_start,
--      ap_idle  => open,
--      ap_ready => open,
--      ap_done  => MatchCalculator_done,
--      bx_V          => bx_out_MatchEngine,
--      bx_o_V        => bx_out_MatchCalculator,
--      bx_o_V_ap_vld => bx_out_MatchCalculator_vld,
--      match_0_dataarray_data_V_ce0         => CM_L3PHIC17_dataarray_data_V_enb,
--      match_0_dataarray_data_V_address0     => CM_L3PHIC17_dataarray_data_V_readaddr,
--      match_0_dataarray_data_V_q0            => CM_L3PHIC17_dataarray_data_V_dout,
--      match_0_nentries_0_V        => CM_L3PHIC17_nentries_0_V_dout(6 downto 0),
--      match_0_nentries_1_V        => CM_L3PHIC17_nentries_1_V_dout(6 downto 0),
--      match_1_dataarray_data_V_ce0         => CM_L3PHIC18_dataarray_data_V_enb,
--      match_1_dataarray_data_V_address0     => CM_L3PHIC18_dataarray_data_V_readaddr,
--      match_1_dataarray_data_V_q0            => CM_L3PHIC18_dataarray_data_V_dout,
--      match_1_nentries_0_V        => CM_L3PHIC18_nentries_0_V_dout(6 downto 0),
--      match_1_nentries_1_V        => CM_L3PHIC18_nentries_1_V_dout(6 downto 0),
--      match_2_dataarray_data_V_ce0         => CM_L3PHIC19_dataarray_data_V_enb,
--      match_2_dataarray_data_V_address0     => CM_L3PHIC19_dataarray_data_V_readaddr,
--      match_2_dataarray_data_V_q0            => CM_L3PHIC19_dataarray_data_V_dout,
--      match_2_nentries_0_V        => CM_L3PHIC19_nentries_0_V_dout(6 downto 0),
--      match_2_nentries_1_V        => CM_L3PHIC19_nentries_1_V_dout(6 downto 0),
--      match_3_dataarray_data_V_ce0         => CM_L3PHIC20_dataarray_data_V_enb,
--      match_3_dataarray_data_V_address0     => CM_L3PHIC20_dataarray_data_V_readaddr,
--      match_3_dataarray_data_V_q0            => CM_L3PHIC20_dataarray_data_V_dout,
--      match_3_nentries_0_V        => CM_L3PHIC20_nentries_0_V_dout(6 downto 0),
--      match_3_nentries_1_V        => CM_L3PHIC20_nentries_1_V_dout(6 downto 0),
--      match_4_dataarray_data_V_ce0         => CM_L3PHIC21_dataarray_data_V_enb,
--      match_4_dataarray_data_V_address0     => CM_L3PHIC21_dataarray_data_V_readaddr,
--      match_4_dataarray_data_V_q0            => CM_L3PHIC21_dataarray_data_V_dout,
--      match_4_nentries_0_V        => CM_L3PHIC21_nentries_0_V_dout(6 downto 0),
--      match_4_nentries_1_V        => CM_L3PHIC21_nentries_1_V_dout(6 downto 0),
--      match_5_dataarray_data_V_ce0         => CM_L3PHIC22_dataarray_data_V_enb,
--      match_5_dataarray_data_V_address0     => CM_L3PHIC22_dataarray_data_V_readaddr,
--      match_5_dataarray_data_V_q0            => CM_L3PHIC22_dataarray_data_V_dout,
--      match_5_nentries_0_V        => CM_L3PHIC22_nentries_0_V_dout(6 downto 0),
--      match_5_nentries_1_V        => CM_L3PHIC22_nentries_1_V_dout(6 downto 0),
--      match_6_dataarray_data_V_ce0         => CM_L3PHIC23_dataarray_data_V_enb,
--      match_6_dataarray_data_V_address0     => CM_L3PHIC23_dataarray_data_V_readaddr,
--      match_6_dataarray_data_V_q0            => CM_L3PHIC23_dataarray_data_V_dout,
--      match_6_nentries_0_V        => CM_L3PHIC23_nentries_0_V_dout(6 downto 0),
--      match_6_nentries_1_V        => CM_L3PHIC23_nentries_1_V_dout(6 downto 0),
--      match_7_dataarray_data_V_ce0         => CM_L3PHIC24_dataarray_data_V_enb,
--      match_7_dataarray_data_V_address0     => CM_L3PHIC24_dataarray_data_V_readaddr,
--      match_7_dataarray_data_V_q0            => CM_L3PHIC24_dataarray_data_V_dout,
--      match_7_nentries_0_V        => CM_L3PHIC24_nentries_0_V_dout(6 downto 0),
--      match_7_nentries_1_V        => CM_L3PHIC24_nentries_1_V_dout(6 downto 0),
--      allstub_dataarray_data_V_ce0         => AS_L3PHICn6_dataarray_data_V_enb,
--      allstub_dataarray_data_V_address0     => AS_L3PHICn6_dataarray_data_V_readaddr,
--      allstub_dataarray_data_V_q0            => AS_L3PHICn6_dataarray_data_V_dout,
--      allproj_dataarray_data_V_ce0         => AP_L3PHIC_dataarray_data_V_enb,
--      allproj_dataarray_data_V_address0     => AP_L3PHIC_dataarray_data_V_readaddr,
--      allproj_dataarray_data_V_q0            => AP_L3PHIC_dataarray_data_V_dout,
--      fullmatch_0_dataarray_data_V_address0 => FM_L1L2_L3PHIC_dataarray_data_V_writeaddr,
--      fullmatch_0_dataarray_data_V_ce0      => open,
--      fullmatch_0_dataarray_data_V_we0      => FM_L1L2_L3PHIC_dataarray_data_V_wea,
--      fullmatch_0_dataarray_data_V_d0       => FM_L1L2_L3PHIC_dataarray_data_V_din,
--      fullmatch_3_dataarray_data_V_address0 => FM_L5L6_L3PHIC_dataarray_data_V_writeaddr,
--      fullmatch_3_dataarray_data_V_ce0      => open,
--      fullmatch_3_dataarray_data_V_we0      => FM_L5L6_L3PHIC_dataarray_data_V_wea,
--      fullmatch_3_dataarray_data_V_d0       => FM_L5L6_L3PHIC_dataarray_data_V_din  );


end rtl;
