--! Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--! User packages
use work.tf_pkg.all;

package memUtil_pkg is

  -- ########################### Types ###########################

  type enum_DL_39 is (negPS10G_2_A,neg2S_3_A,negPS_1_A,PS10G_2_A,neg2S_4_B,negPS_2_A,twoS_2_B,twoS_4_B,PS10G_3_A,twoS_2_A,PS10G_1_A,PS_1_A,neg2S_4_A,twoS_1_B,negPS10G_1_A,PS_1_B,twoS_3_B,PS10G_2_B,negPS10G_3_A,PS10G_1_B,neg2S_1_B,neg2S_1_A,negPS_1_B,neg2S_2_B,PS10G_3_B,PS_2_A,neg2S_3_B,twoS_1_A,negPS10G_3_B,negPS10G_2_B,PS_2_B,neg2S_2_A,negPS_2_B,negPS10G_1_B,twoS_3_A,twoS_4_A);

  type enum_IL_36 is (L1PHIH_PS10G_2_B,L3PHIB_negPS_2_B,L6PHIB_neg2S_4_A,L1PHID_PS10G_1_A,L6PHIC_neg2S_3_B,L6PHIC_neg2S_4_B,L2PHIC_PS10G_3_A,L1PHIH_negPS10G_2_B,L1PHID_PS10G_2_A,L3PHIA_negPS_1_A,L5PHID_2S_2_B,L5PHIC_neg2S_1_B,L2PHIB_negPS10G_3_A,L6PHIB_2S_3_B,L1PHIF_negPS10G_2_B,L5PHIC_neg2S_2_B,L4PHIC_neg2S_1_B,L3PHID_PS_2_B,L6PHIC_2S_3_B,L2PHIB_PS10G_3_A,L3PHIA_PS_1_A,L6PHIB_neg2S_3_A,L5PHIB_neg2S_2_B,L6PHIB_2S_4_A,L5PHIC_2S_2_A,L1PHIF_PS10G_1_B,L2PHIA_PS10G_3_A,L1PHIC_negPS10G_2_B,L6PHIA_2S_3_A,L1PHIE_PS10G_2_A,L1PHIA_negPS10G_1_A,L1PHIB_negPS10G_1_A,L6PHIB_2S_3_A,L1PHIF_PS10G_2_A,L3PHIB_PS_1_A,L1PHIH_negPS10G_1_B,L1PHIE_PS10G_2_B,L5PHIB_neg2S_2_A,L5PHIB_neg2S_1_A,L4PHIA_2S_1_A,L6PHIC_2S_3_A,L1PHIF_PS10G_1_A,L5PHIB_2S_2_A,L3PHID_PS_1_B,L1PHIG_PS10G_2_B,L3PHIC_negPS_2_A,L1PHIA_PS10G_1_A,L1PHIC_negPS10G_1_A,L2PHIB_PS10G_3_B,L3PHID_negPS_2_B,L1PHIB_PS10G_2_A,L5PHID_neg2S_1_B,L4PHIC_2S_1_B,L1PHIE_negPS10G_1_B,L2PHIA_negPS10G_3_A,L1PHID_negPS10G_2_B,L5PHIC_2S_1_B,L3PHIB_negPS_1_A,L5PHIA_neg2S_1_A,L3PHID_negPS_1_B,L4PHID_2S_1_B,L1PHIC_negPS10G_1_B,L1PHID_negPS10G_1_B,L1PHIG_PS10G_1_A,L2PHIB_negPS10G_3_B,L1PHID_PS10G_2_B,L1PHIE_PS10G_1_B,L4PHIB_neg2S_1_B,L1PHIF_negPS10G_2_A,L5PHID_2S_1_B,L1PHIG_PS10G_1_B,L3PHIB_PS_2_A,L1PHIC_PS10G_1_A,L3PHIC_PS_2_A,L1PHIG_negPS10G_2_B,L1PHIF_negPS10G_1_B,L6PHIA_2S_4_A,L5PHIC_2S_2_B,L2PHID_PS10G_3_B,L3PHIB_negPS_2_A,L6PHID_2S_4_B,L1PHIE_negPS10G_2_B,L1PHIB_PS10G_1_A,L4PHID_neg2S_1_B,L1PHIC_PS10G_2_B,L1PHIC_negPS10G_2_A,L5PHIA_neg2S_2_A,L4PHIB_neg2S_1_A,L3PHIB_PS_1_B,L1PHIB_negPS10G_2_A,L1PHIH_PS10G_1_B,L4PHIC_2S_1_A,L6PHIB_neg2S_3_B,L3PHIC_PS_2_B,L3PHIB_PS_2_B,L6PHID_neg2S_4_B,L3PHIA_PS_2_A,L5PHIB_2S_1_A,L1PHIF_PS10G_2_B,L5PHIA_2S_1_A,L3PHIC_PS_1_B,L4PHIC_neg2S_1_A,L1PHIA_PS10G_2_A,L6PHIB_neg2S_4_B,L1PHID_negPS10G_2_A,L4PHIB_2S_1_B,L1PHIA_negPS10G_2_A,L6PHID_neg2S_3_B,L6PHIC_2S_4_B,L2PHIC_negPS10G_3_A,L6PHIC_neg2S_3_A,L2PHID_negPS10G_3_B,L3PHIC_negPS_1_B,L3PHIB_negPS_1_B,L3PHIA_negPS_2_A,L5PHID_neg2S_2_B,L5PHIB_2S_2_B,L5PHIC_neg2S_2_A,L1PHIE_negPS10G_2_A,L6PHIB_2S_4_B,L4PHIB_2S_1_A,L3PHIC_negPS_2_B,L6PHIC_2S_4_A,L3PHIC_PS_1_A,L2PHIC_negPS10G_3_B,L6PHID_2S_3_B,L4PHIA_neg2S_1_A,L1PHIC_PS10G_2_A,L1PHIG_negPS10G_1_B,L6PHIA_neg2S_4_A,L1PHIE_PS10G_1_A,L6PHIC_neg2S_4_A,L2PHIC_PS10G_3_B,L5PHIA_2S_2_A,L1PHID_negPS10G_1_A,L6PHIA_neg2S_3_A);

  type enum_AS_36 is (L4PHIDn2,L3PHICn6,L5PHIBn1,L3PHIDn1,L1PHIHn3,L1PHIBn1,L1PHIAn1,L2PHICn6,L1PHIGn3,L4PHIAn3,L2PHICn4,L2PHICn2,L1PHIDn2,L3PHICn2,L4PHIBn4,L2PHIDn4,L4PHIBn1,L5PHIAn2,L1PHIDn1,L4PHIDn1,L1PHICn3,L1PHICn4,L1PHIGn2,L2PHIBn3,L3PHIBn2,L3PHICn4,L1PHIEn1,L6PHIDn3,L1PHIFn3,L1PHIAn3,L2PHICn7,L6PHICn2,L2PHIBn6,L5PHIBn3,L2PHICn1,L3PHIDn3,L4PHICn4,L1PHIBn2,L4PHIAn2,L2PHIBn1,L5PHIDn2,L2PHIAn6,L3PHIDn2,L2PHIBn7,L3PHIBn6,L2PHICn5,L2PHIAn1,L2PHIBn8,L2PHIBn5,L6PHIBn3,L1PHIFn1,L6PHIAn2,L6PHIDn2,L5PHICn1,L5PHIDn1,L1PHIHn2,L1PHIEn3,L4PHIBn3,L4PHIAn1,L5PHICn3,L4PHIBn2,L3PHIBn5,L3PHIBn4,L3PHICn3,L1PHIFn4,L6PHICn1,L2PHIAn5,L3PHIBn3,L3PHICn1,L2PHIBn2,L5PHIBn2,L6PHIBn2,L4PHIDn3,L1PHICn2,L6PHICn3,L6PHICn4,L2PHICn3,L1PHIFn2,L4PHICn3,L2PHIDn2,L3PHIDn4,L1PHIGn1,L6PHIDn1,L2PHIAn3,L6PHIBn1,L1PHIHn1,L2PHIAn4,L2PHIDn3,L3PHIAn2,L1PHIAn2,L3PHIBn1,L2PHIDn1,L5PHIAn1,L2PHIAn2,L6PHIAn3,L1PHICn1,L2PHIBn4,L4PHICn2,L6PHIBn4,L3PHIAn3,L1PHIDn3,L1PHIBn3,L4PHICn1,L6PHIAn1,L2PHIDn6,L3PHICn5,L2PHIDn5,L5PHICn2,L3PHIAn1,L1PHIEn2);

  type enum_VMSME_17 is (L5PHID28n1,L5PHIC23n1,L4PHIB15n1,L4PHIC21n1,L4PHIA4n1,L5PHID25n1,L6PHIB12n1,L6PHIC18n1,L4PHIB14n1,L4PHIA3n1,L4PHIB10n1,L5PHIB13n1,L6PHIB9n1,L6PHID32n1,L5PHIA5n1,L5PHIA1n1,L4PHID28n1,L5PHIC17n1,L4PHID25n1,L4PHIC22n1,L6PHIA2n1,L6PHIA6n1,L4PHIA7n1,L6PHIC21n1,L5PHIC22n1,L4PHIB9n1,L4PHID30n1,L5PHIB14n1,L6PHIB16n1,L6PHID26n1,L6PHIA3n1,L6PHIC17n1,L5PHID31n1,L6PHIC22n1,L6PHID30n1,L6PHID31n1,L5PHIB15n1,L4PHIC24n1,L5PHID32n1,L4PHIC17n1,L4PHID29n1,L4PHIA6n1,L4PHID27n1,L6PHIB13n1,L6PHIC24n1,L5PHIB11n1,L5PHID26n1,L4PHIC20n1,L5PHIC24n1,L5PHIA2n1,L5PHID30n1,L5PHIB10n1,L6PHIC19n1,L5PHIA6n1,L4PHID31n1,L5PHID29n1,L5PHIA8n1,L4PHIA8n1,L4PHIB16n1,L4PHID32n1,L6PHIB11n1,L5PHIC20n1,L4PHID26n1,L4PHIB13n1,L6PHIC23n1,L6PHIA8n1,L4PHIA2n1,L5PHID27n1,L6PHIA4n1,L5PHIB16n1,L5PHIC21n1,L5PHIC19n1,L6PHIB10n1,L6PHIB15n1,L6PHIB14n1,L5PHIA3n1,L5PHIA4n1,L5PHIB12n1,L4PHIB11n1,L6PHID28n1,L4PHIB12n1,L5PHIC18n1,L4PHIC19n1,L6PHIA7n1,L4PHIA1n1,L6PHIA5n1,L6PHID29n1,L4PHIC18n1,L5PHIB9n1,L4PHIC23n1,L6PHID27n1,L6PHID25n1,L6PHIC20n1,L5PHIA7n1,L4PHIA5n1,L6PHIA1n1);

  type enum_VMSME_16 is (L2PHIC21n1,L2PHID31n1,L2PHIB10n1,L1PHIF22n1,L3PHID25n1,L1PHIA2n1,L1PHID15n1,L1PHIA3n1,L3PHIA3n1,L3PHIC23n1,L1PHID16n1,L1PHIE17n1,L3PHID26n1,L2PHID29n1,L2PHID30n1,L2PHIA4n1,L1PHIG28n1,L2PHIC19n1,L1PHIA4n1,L1PHIC9n1,L3PHIB11n1,L1PHIF21n1,L1PHIF23n1,L1PHIE19n1,L2PHIC24n1,L2PHIB9n1,L3PHIC21n1,L3PHIA5n1,L3PHIB10n1,L3PHID28n1,L3PHID32n1,L3PHID30n1,L2PHIB14n1,L2PHIC17n1,L1PHIH30n1,L1PHIG25n1,L1PHIH31n1,L3PHIA4n1,L3PHIA7n1,L2PHIB16n1,L3PHIC17n1,L1PHIH32n1,L2PHIC18n1,L2PHIA7n1,L3PHIA6n1,L3PHIA8n1,L3PHIB9n1,L2PHID32n1,L3PHIC22n1,L1PHIC10n1,L2PHIA5n1,L2PHIC23n1,L1PHIA1n1,L1PHIC12n1,L1PHIC11n1,L1PHID13n1,L2PHIC20n1,L2PHIA6n1,L3PHIC18n1,L1PHIE20n1,L2PHIA3n1,L3PHIB14n1,L2PHIA8n1,L1PHIB7n1,L1PHIB5n1,L1PHIB8n1,L2PHID26n1,L1PHIG26n1,L2PHIB13n1,L2PHIB15n1,L2PHID28n1,L3PHID29n1,L1PHID14n1,L1PHIB6n1,L2PHIA2n1,L3PHIB15n1,L3PHID31n1,L3PHIC24n1,L2PHIA1n1,L3PHIA1n1,L3PHIC19n1,L1PHIE18n1,L1PHIG27n1,L3PHIB16n1,L3PHIB13n1,L2PHIB11n1,L2PHIB12n1,L1PHIH29n1,L2PHID25n1,L2PHID27n1,L1PHIF24n1,L3PHID27n1,L3PHIB12n1,L3PHIC20n1,L2PHIC22n1,L3PHIA2n1);

  type enum_VMSTE_22 is (L2PHIJ6n3,L3PHID15n2,L2PHIJ6n2,L3PHID13n5,L1PHIA2n3,L1PHIB6n2,L1PHIB8n3,L1PHIA4n2,L3PHID14n3,L1PHIE19n3,L2PHIK10n2,L1PHIB6n3,L1PHIE17n4,L1PHID16n3,L3PHIC9n5,L1PHIG25n3,L3PHID16n3,L1PHID16n4,L2PHIK12n1,L1PHIA1n3,L1PHIF23n2,L1PHIH31n4,L1PHIC12n1,L1PHIG25n2,L1PHIG26n3,L1PHIB7n1,L3PHIA2n4,L3PHIA2n5,L2PHII3n3,L1PHIF21n4,L1PHIB8n2,L3PHIA3n1,L1PHIH32n2,L3PHIC10n6,L3PHIC11n6,L2PHIL13n1,L2PHIL15n3,L3PHIB5n3,L2PHIJ8n1,L1PHIH32n3,L1PHIF24n2,L1PHIA1n2,L1PHIF23n5,L2PHIJ8n3,L1PHIG27n2,L1PHIG26n2,L1PHIA4n1,L3PHID16n2,L1PHIB6n5,L3PHIA1n4,L2PHIL16n1,L1PHIG28n2,L2PHIL13n3,L3PHIA4n1,L3PHID14n5,L1PHIG27n4,L2PHIK12n2,L1PHIC11n4,L3PHIC11n5,L3PHIB6n2,L1PHIB5n2,L3PHIC9n6,L1PHIC11n1,L1PHIF22n1,L1PHIC11n2,L3PHID15n1,L1PHIG27n5,L3PHID15n3,L1PHIE17n3,L1PHIC12n3,L1PHIB5n1,L1PHIC10n4,L1PHID14n2,L1PHIC9n3,L3PHIB6n5,L1PHIH29n1,L1PHID14n4,L1PHIE17n5,L1PHIB8n1,L1PHIE20n4,L1PHIG28n1,L3PHIC12n4,L1PHIA3n4,L1PHID15n1,L1PHIE17n1,L3PHIB5n5,L1PHIG25n4,L3PHID16n4,L1PHIE20n3,L1PHID16n2,L3PHIC12n5,L2PHIK11n2,L3PHID13n3,L3PHIB7n2,L1PHIF23n4,L1PHIC10n5,L3PHID13n2,L2PHII4n1,L3PHIB6n4,L2PHII3n1,L2PHII1n2,L2PHIL14n1,L1PHIA4n4,L1PHIE18n1,L3PHIA3n2,L2PHIK9n3,L3PHIC11n1,L2PHII3n2,L1PHIE18n2,L1PHIH32n1,L1PHID13n2,L3PHIC10n3,L1PHIH30n4,L1PHIA3n2,L1PHIE17n2,L1PHIB6n1,L3PHID14n4,L2PHIK10n1,L1PHIF24n5,L2PHII4n3,L2PHIK9n1,L2PHIJ7n2,L3PHIB7n4,L3PHID13n1,L3PHIC12n3,L1PHIC10n1,L3PHIB8n2,L2PHIJ5n1,L2PHIJ6n1,L1PHIF21n1,L1PHIF21n3,L1PHIC9n5,L1PHIF22n2,L1PHIC12n2,L1PHIH31n1,L1PHIG25n5,L1PHIB7n4,L1PHIA4n3,L3PHIB5n4,L1PHID13n1,L1PHIF24n3,L1PHIG28n5,L1PHIE18n4,L3PHIB7n3,L2PHIL14n2,L2PHIK11n3,L3PHIC9n2,L3PHIC11n3,L3PHIB7n1,L1PHIE19n2,L3PHIA4n3,L1PHID13n4,L1PHIF24n4,L2PHIK12n3,L3PHIB8n4,L3PHIB7n6,L1PHIH30n5,L2PHIJ8n2,L1PHIC11n3,L1PHIH30n1,L3PHIC10n5,L3PHID15n6,L1PHIC10n2,L1PHIC10n3,L3PHID16n1,L1PHIG28n4,L1PHID13n5,L1PHIG28n3,L3PHIC9n1,L1PHID15n5,L1PHIH29n2,L3PHIA3n3,L1PHIH30n3,L3PHIA3n4,L1PHIA4n5,L1PHIF22n3,L1PHID14n5,L3PHIA3n5,L1PHIA3n5,L1PHIH31n3,L2PHIJ5n2,L1PHIB7n5,L2PHIL15n1,L1PHIA3n1,L1PHIF22n5,L2PHIL14n3,L2PHII2n1,L1PHID15n3,L1PHIG27n1,L3PHIC12n2,L1PHIC12n4,L3PHIA2n1,L1PHIB5n3,L3PHIA1n2,L3PHIC11n4,L1PHIF23n3,L1PHIH30n2,L1PHIF21n5,L1PHIA2n4,L3PHIC12n6,L3PHIB5n2,L3PHIA1n3,L1PHIH29n5,L1PHIB5n5,L3PHIB7n5,L3PHIA4n6,L1PHIF21n2,L3PHIA2n2,L1PHIH31n2,L1PHIF24n1,L1PHIC9n2,L3PHIC9n4,L3PHIA1n1,L3PHID13n6,L3PHIC12n1,L1PHIA2n1,L1PHIB8n5,L3PHIA3n6,L3PHID14n2,L1PHIC12n5,L2PHII1n1,L2PHIJ5n3,L1PHIB6n4,L3PHIB5n6,L3PHIC11n2,L1PHIF22n4,L2PHII2n2,L2PHIL16n2,L1PHIB7n2,L2PHIK9n2,L3PHIA4n4,L2PHIL13n2,L3PHIC10n2,L3PHIB8n1,L1PHIA3n3,L3PHIC10n1,L3PHID15n4,L1PHIE20n5,L1PHID13n3,L1PHIE18n5,L2PHIL15n2,L1PHIE20n1,L1PHID16n5,L3PHID15n5,L3PHIB6n3,L3PHID14n6,L1PHIB7n3,L3PHIB6n6,L1PHIA1n1,L1PHIE19n4,L1PHIH29n3,L1PHID14n3,L1PHIE19n1,L1PHIB8n4,L3PHID14n1,L1PHIG26n4,L1PHIE19n5,L1PHIA2n2,L2PHIK11n1,L3PHIC10n4,L1PHID16n1,L3PHIA2n3,L3PHIB8n6,L1PHIC11n5,L1PHIE20n2,L3PHIA4n2,L1PHID14n1,L2PHII2n3,L3PHIB5n1,L2PHIK10n3,L1PHIE18n3,L1PHIC9n1,L3PHID13n4,L3PHIA2n6,L2PHIJ7n3,L2PHIJ7n1,L1PHIC9n4,L1PHIG26n1,L3PHIB6n1,L1PHIG27n3,L1PHID15n2,L1PHIG26n5,L1PHID15n4,L3PHIB8n5,L1PHIF23n1,L3PHIB8n3,L2PHII4n2,L3PHIA4n5,L1PHIG25n1,L1PHIB5n4,L1PHIH29n4,L3PHIC9n3);

  type enum_VMSTE_17 is (L6PHIC22n1,L6PHID27n1,L6PHID26n1,L6PHIC24n2,L6PHIB11n4,L6PHIA6n3,L6PHIB13n2,L6PHIA8n3,L6PHID25n1,L6PHIB15n3,L6PHID29n1,L6PHIB14n3,L4PHID25n2,L6PHIB12n1,L4PHIA4n1,L6PHIB15n1,L4PHIA6n1,L6PHID25n3,L6PHID27n4,L6PHIC17n3,L4PHIC18n1,L6PHID25n2,L6PHIB12n4,L6PHID28n1,L6PHIC19n1,L4PHIC22n2,L6PHID29n4,L6PHIC19n2,L6PHIB14n2,L6PHIB11n1,L6PHIC18n1,L6PHIB9n2,L4PHIC20n2,L6PHIB10n3,L4PHIC18n3,L4PHIB13n3,L4PHIB14n3,L4PHIB14n2,L4PHIB13n2,L4PHIB16n2,L6PHIA3n3,L4PHIC17n3,L6PHID27n2,L6PHIB11n3,L6PHIB12n2,L6PHID28n2,L6PHIA7n3,L4PHID25n1,L4PHIC20n1,L4PHID32n2,L4PHIB9n1,L4PHIA7n3,L6PHIB14n1,L4PHID30n2,L4PHIA4n2,L6PHIA6n1,L4PHID29n1,L4PHIA6n3,L6PHID31n1,L6PHIA4n3,L6PHIC18n4,L6PHID29n3,L6PHIC17n2,L4PHID27n3,L4PHIC20n3,L4PHIC19n2,L4PHIB10n3,L4PHIC19n3,L6PHIA1n2,L6PHIA7n2,L6PHIC23n1,L4PHIB15n3,L6PHIB16n2,L6PHIC20n1,L4PHIC17n2,L4PHIB12n3,L6PHIA8n4,L6PHIC23n2,L4PHIC21n3,L4PHIB10n1,L6PHIA7n1,L6PHIC20n3,L4PHIB15n1,L6PHID26n3,L6PHIC22n2,L4PHID28n3,L6PHIA5n1,L6PHID32n1,L4PHID26n3,L6PHIB11n2,L6PHIA4n1,L4PHID30n3,L4PHID29n2,L6PHIC23n3,L6PHIC18n3,L6PHIA8n2,L6PHIA3n2,L4PHID26n2,L4PHID28n2,L4PHID31n2,L6PHIB16n1,L6PHID31n3,L6PHIC18n2,L4PHIB9n2,L4PHIA8n1,L4PHIC23n1,L6PHID27n3,L4PHID32n1,L4PHIB11n1,L6PHID26n4,L6PHID31n2,L6PHIA2n2,L6PHIC21n3,L4PHIB12n1,L6PHID32n2,L6PHID25n4,L6PHIA2n1,L4PHIA5n3,L6PHID28n4,L4PHIC23n2,L4PHIB12n2,L6PHIB10n1,L4PHIC21n2,L6PHIB10n2,L4PHIC24n1,L6PHIA6n2,L6PHIC22n3,L6PHIB13n1,L4PHIB9n3,L4PHIB16n1,L6PHID30n1,L4PHID29n3,L6PHIA6n4,L6PHIB15n2,L4PHID30n1,L6PHIC20n4,L6PHIC22n4,L6PHIB15n4,L4PHIB16n3,L4PHIC19n1,L4PHIA2n1,L6PHIC19n4,L6PHIC21n2,L6PHIC21n1,L4PHIB14n1,L6PHIB16n4,L4PHIA6n2,L4PHID26n1,L6PHIC24n1,L4PHIA8n2,L6PHIA3n1,L6PHIA4n4,L6PHIB9n3,L6PHIB10n4,L4PHIB13n1,L4PHID25n3,L6PHIA2n3,L6PHID29n2,L4PHIC22n1,L6PHIC20n2,L4PHIC23n3,L6PHIC23n4,L4PHIA3n3,L4PHIC17n1,L6PHIB13n3,L4PHIA4n3,L4PHIA3n1,L6PHID30n2,L4PHIA8n3,L4PHIA7n2,L6PHIC17n1,L4PHIA1n1,L4PHID27n2,L4PHIA1n2,L6PHIA5n3,L6PHID26n2,L6PHIC24n3,L4PHIA2n2,L6PHID30n3,L4PHIC24n3,L4PHID28n1,L6PHIB14n4,L6PHIB9n1,L6PHIC24n4,L6PHIA1n1,L4PHIB15n2,L6PHIB16n3,L6PHIA5n4,L4PHID31n1,L4PHIA5n2,L6PHIA5n2,L6PHIB13n4,L4PHIB11n2,L4PHID27n1,L4PHIA3n2,L4PHIC21n1,L6PHIA4n2,L4PHIA7n1,L6PHIC17n4,L4PHIC18n2,L4PHIB11n3,L6PHIB12n3,L6PHIC21n4,L4PHIC24n2,L4PHIA5n1,L6PHIB9n4,L4PHIB10n2,L4PHIC22n3,L6PHIA8n1,L6PHID28n3,L6PHIC19n3,L6PHIA7n4);

  type enum_VMSTE_23 is (L5PHIB7n1,L5PHIC10n3,L5PHID15n1,L5PHIB6n4,L5PHIB8n8,L5PHIC12n6,L5PHID16n5,L5PHIC11n5,L5PHID15n3,L5PHIA3n7,L5PHID14n2,L5PHID13n5,L5PHIA4n8,L5PHIB8n7,L5PHIA3n5,L5PHIB5n3,L5PHIC12n2,L5PHIB8n4,L5PHIC9n1,L5PHIC10n8,L5PHID16n2,L5PHIC12n5,L5PHIB6n2,L5PHIC9n4,L5PHIA1n1,L5PHIB7n8,L5PHIA4n4,L5PHIB7n4,L5PHID13n3,L5PHIB6n1,L5PHID15n4,L5PHIC11n1,L5PHIA4n6,L5PHIC12n4,L5PHIC11n2,L5PHIA3n4,L5PHID13n4,L5PHID13n2,L5PHIB5n8,L5PHIC9n3,L5PHIA3n6,L5PHID14n5,L5PHIC11n8,L5PHIA2n6,L5PHIB8n3,L5PHIC11n4,L5PHIC12n1,L5PHIA1n2,L5PHIB7n2,L5PHIA2n7,L5PHIA3n2,L5PHIA4n2,L5PHIB5n2,L5PHIA3n8,L5PHIC11n6,L5PHID14n4,L5PHIA2n2,L5PHID16n1,L5PHID13n7,L5PHIA2n5,L5PHID14n7,L5PHIC12n8,L5PHIA2n4,L5PHID13n1,L5PHIB7n5,L5PHIC10n7,L5PHIA1n4,L5PHIC9n6,L5PHID16n4,L5PHIA2n1,L5PHIC10n2,L5PHIA4n3,L5PHIC12n3,L5PHIB7n3,L5PHIB6n8,L5PHIB8n1,L5PHIB6n3,L5PHIA2n3,L5PHIC12n7,L5PHIC11n7,L5PHIC9n5,L5PHIC9n7,L5PHID13n8,L5PHIC11n3,L5PHIC9n2,L5PHIC10n1,L5PHIB5n6,L5PHIC10n5,L5PHIB5n1,L5PHIA3n1,L5PHIA4n7,L5PHID14n3,L5PHIC10n4,L5PHIB8n2,L5PHIA1n5,L5PHIB5n5,L5PHID15n7,L5PHIA3n3,L5PHID16n3,L5PHID14n1,L5PHIB5n7,L5PHIB6n6,L5PHIA4n1,L5PHIB8n6,L5PHID14n6,L5PHID15n2,L5PHIA4n5,L5PHIB6n5,L5PHID15n6,L5PHIB7n7,L5PHID15n5,L5PHIC9n8,L5PHID14n8,L5PHID13n6,L5PHIB7n6,L5PHIC10n6,L5PHIB8n5,L5PHIA1n3,L5PHIB5n4,L5PHIB6n7);

  type enum_VMSTE_16 is (L2PHID28n3,L2PHID30n1,L2PHID27n2,L2PHIC23n3,L2PHIB13n3,L3PHIJ7n3,L2PHIA8n4,L3PHIJ8n1,L2PHIB9n5,L2PHIC20n5,L2PHIC22n1,L2PHIB10n1,L3PHII1n1,L2PHIB12n3,L2PHIB9n4,L3PHIK9n3,L2PHIC22n2,L2PHID32n2,L2PHIC24n1,L2PHID30n4,L3PHII3n3,L3PHII1n2,L2PHID30n2,L3PHIK11n2,L2PHIC22n4,L2PHIA2n2,L3PHIL14n3,L2PHIB16n3,L2PHID30n3,L2PHIA4n2,L2PHID28n2,L3PHIK10n2,L2PHIC18n1,L2PHIB15n1,L2PHIC22n3,L2PHIC22n5,L2PHID32n3,L2PHIB14n4,L2PHIA4n3,L2PHIB16n2,L3PHIJ8n3,L2PHIB16n4,L2PHIB15n4,L2PHIA3n3,L2PHIB10n2,L3PHIJ5n3,L2PHIB12n1,L2PHIC21n2,L2PHID27n3,L2PHIA5n1,L2PHIB12n5,L2PHID25n2,L2PHIC23n5,L2PHIB11n3,L3PHIJ6n3,L2PHIC17n4,L2PHIB10n5,L3PHIL15n1,L2PHIA8n3,L3PHIK9n2,L3PHII4n3,L2PHIA4n1,L2PHIA7n5,L2PHID27n4,L2PHIA1n1,L2PHID29n1,L2PHIC23n1,L2PHIA2n1,L2PHIC19n2,L2PHID29n2,L2PHIC23n4,L2PHID26n3,L2PHIA3n1,L2PHIB11n4,L2PHIC18n5,L3PHIL15n3,L2PHID25n3,L2PHIC17n1,L2PHID28n4,L2PHIC17n2,L2PHIC24n5,L2PHIC19n1,L2PHIB12n4,L2PHIC24n3,L3PHII2n1,L2PHIA1n2,L2PHID28n1,L2PHIB13n2,L2PHID26n1,L2PHIC20n2,L3PHIL13n2,L2PHID26n5,L2PHIA5n3,L2PHIB10n4,L2PHIA8n5,L3PHIJ7n1,L2PHIA7n4,L2PHID27n5,L3PHII3n1,L2PHIC18n2,L2PHIA3n2,L3PHIK11n3,L2PHIA5n4,L2PHIA4n4,L2PHIC21n3,L2PHIA2n4,L3PHIK10n3,L2PHIC19n4,L2PHIB11n1,L2PHIA6n3,L2PHIB14n5,L2PHIB9n1,L3PHIK12n3,L2PHIB15n3,L2PHID32n1,L2PHIC19n3,L3PHIJ8n2,L3PHIK12n2,L2PHIA5n5,L2PHIA1n3,L2PHIB14n2,L2PHIC21n5,L3PHIL15n2,L2PHID26n2,L2PHIA6n2,L3PHII3n2,L2PHIB10n3,L2PHIB13n5,L3PHII2n2,L3PHIJ7n2,L2PHIC20n3,L3PHII4n1,L2PHID26n4,L2PHIA7n1,L2PHIA8n2,L2PHIB11n2,L2PHIC21n1,L2PHID31n3,L2PHIC17n3,L2PHID27n1,L2PHID29n5,L2PHID31n2,L2PHIB9n3,L2PHIB15n2,L2PHIC18n3,L3PHIL13n3,L2PHIA7n2,L2PHIA3n4,L2PHID31n4,L2PHIC20n4,L2PHIC19n5,L2PHIB13n1,L2PHIB12n2,L2PHIB13n4,L3PHIL16n2,L3PHIL14n2,L2PHIA5n2,L3PHIJ6n2,L2PHIC24n4,L2PHIA6n5,L2PHIC17n5,L3PHIL13n1,L3PHIL16n1,L2PHIA8n1,L2PHID25n1,L2PHIA4n5,L2PHIB16n5,L2PHIB14n3,L2PHID28n5,L2PHID25n5,L2PHID29n4,L2PHIB14n1,L2PHIA2n3,L3PHII4n2,L2PHIB11n5,L2PHIB15n5,L2PHIA7n3,L2PHIC18n4,L3PHIL14n1,L2PHID29n3,L2PHID30n5,L3PHIK10n1,L3PHIK11n1,L2PHIA6n4,L2PHID31n1,L3PHIJ5n1,L2PHIA6n1,L2PHIC20n1,L2PHIC23n2,L3PHIJ5n2,L2PHIC24n2,L3PHIJ6n1,L2PHIB16n1,L2PHIB9n2,L2PHID25n4,L2PHIA3n5,L3PHIK9n1,L2PHIC21n4,L3PHII2n3,L3PHIK12n1);

  type enum_SP_14 is (L3PHID14_L4PHID29,L3PHID14_L4PHID25,L1PHIF21_L2PHIC22,L1PHIE18_L2PHIB16,L3PHIC9_L4PHIC17,L5PHIA1_L6PHIA2,L3PHID13_L4PHID26,L2PHII4_L3PHII4,L5PHIC11_L6PHIC23,L2PHIK12_L3PHIK12,L5PHIB6_L6PHIB10,L3PHIA1_L4PHIA3,L3PHIA1_L4PHIA1,L1PHIA2_L2PHIA2,L3PHIB5_L4PHIA8,L3PHIC11_L4PHIC20,L1PHIG26_L2PHID27,L5PHID14_L6PHID26,L1PHIH31_L2PHID29,L1PHIC10_L2PHIB9,L1PHIC12_L2PHIB12,L3PHIB8_L4PHIB14,L3PHIA3_L4PHIA5,L1PHIF23_L2PHID25,L2PHIJ5_L3PHIJ5,L5PHIA3_L6PHIA6,L1PHIE19_L2PHIC17,L3PHIB7_L4PHIB11,L2PHII3_L3PHII3,L5PHIB8_L6PHIC18,L1PHIG25_L2PHID26,L1PHIB7_L2PHIB9,L1PHIA4_L2PHIA6,L3PHIA4_L4PHIA5,L1PHIE17_L2PHIB16,L1PHID15_L2PHIC17,L5PHID13_L6PHID27,L5PHIB8_L6PHIB13,L1PHIF24_L2PHIC24,L1PHIG26_L2PHID28,L3PHIC11_L4PHIC24,L2PHII3_L3PHII2,L1PHIG28_L2PHID30,L5PHIB8_L6PHIB14,L5PHIB6_L6PHIB13,L3PHIA3_L4PHIA3,L1PHIF21_L2PHIC21,L2PHIK10_L3PHIK10,L5PHIB5_L6PHIB12,L5PHIC12_L6PHIC21,L3PHIA3_L4PHIA4,L5PHIC12_L6PHIC24,L3PHIC12_L4PHIC22,L1PHIA1_L2PHIA3,L5PHID16_L6PHID29,L5PHID16_L6PHID32,L3PHIC12_L4PHIC21,L5PHID15_L6PHID29,L3PHIA4_L4PHIA8,L3PHIB5_L4PHIA7,L5PHID14_L6PHID28,L2PHIL15_L3PHIL14,L5PHIC12_L6PHIC23,L3PHIA1_L4PHIA4,L1PHID16_L2PHIB15,L1PHIC10_L2PHIB11,L1PHIF24_L2PHIC22,L3PHIA3_L4PHIA7,L5PHIA4_L6PHIA6,L5PHID13_L6PHID29,L5PHIC12_L6PHIC20,L3PHIA2_L4PHIA2,L1PHIH30_L2PHID30,L5PHIC10_L6PHIC18,L5PHIC11_L6PHIC18,L1PHIE18_L2PHIC20,L3PHIC11_L4PHIC21,L3PHIA4_L4PHIA7,L3PHID13_L4PHID25,L3PHIC12_L4PHIC23,L1PHIC9_L2PHIB9,L5PHIA4_L6PHIA8,L1PHIA4_L2PHIA5,L1PHID16_L2PHIB14,L3PHIB6_L4PHIB10,L5PHID14_L6PHID31,L1PHIH32_L2PHID32,L2PHIL14_L3PHIL15,L3PHIA2_L4PHIA1,L2PHIK12_L3PHIL13,L3PHIC9_L4PHIC19,L3PHIA4_L4PHIA6,L5PHIC12_L6PHID27,L1PHIE19_L2PHIC20,L3PHIC10_L4PHIC21,L1PHIB8_L2PHIB10,L1PHIG28_L2PHID29,L1PHIB5_L2PHIA6,L5PHIC10_L6PHIC20,L1PHIA3_L2PHIA2,L5PHIB6_L6PHIB12,L5PHIB8_L6PHIC19,L2PHII1_L3PHII2,L5PHIB8_L6PHIB12,L5PHIA3_L6PHIA5,L1PHIG27_L2PHID28,L1PHIC12_L2PHIB11,L5PHID15_L6PHID27,L1PHIF24_L2PHIC23,L1PHIB8_L2PHIA6,L1PHIG25_L2PHID27,L2PHII4_L3PHII3,L1PHIC9_L2PHIA7,L3PHID15_L4PHID32,L1PHIA4_L2PHIA4,L1PHIA3_L2PHIA4,L3PHID16_L4PHID30,L1PHIG27_L2PHID29,L5PHID16_L6PHID28,L5PHIA4_L6PHIA4,L3PHIC10_L4PHIC20,L3PHIC10_L4PHIC18,L1PHIH32_L2PHID30,L1PHIF22_L2PHIC23,L5PHIC11_L6PHIC20,L1PHIC9_L2PHIB11,L1PHIF23_L2PHIC24,L5PHID13_L6PHIC23,L1PHID13_L2PHIB13,L5PHID14_L6PHIC24,L1PHIF21_L2PHIC23,L1PHIG28_L2PHID27,L1PHIE17_L2PHIB15,L1PHIE18_L2PHIC17,L5PHIB6_L6PHIB9,L5PHIB8_L6PHIB16,L1PHIF23_L2PHIC23,L1PHIB5_L2PHIA7,L1PHIH29_L2PHID28,L5PHIC12_L6PHIC22,L2PHIK11_L3PHIK10,L5PHID13_L6PHID26,L5PHID15_L6PHID28,L1PHID14_L2PHIB14,L2PHII2_L3PHII2,L2PHIK11_L3PHIK11,L1PHID15_L2PHIB14,L5PHIC10_L6PHIC23,L5PHIC11_L6PHID25,L1PHIA1_L2PHIA2,L5PHID13_L6PHIC24,L1PHID13_L2PHIB12,L3PHIC9_L4PHIC18,L5PHID15_L6PHID31,L1PHIE18_L2PHIC18,L5PHIB8_L6PHIC17,L1PHIE18_L2PHIC19,L1PHIC11_L2PHIB12,L2PHII3_L3PHII4,L5PHIC9_L6PHIC21,L1PHIG25_L2PHID25,L1PHIB7_L2PHIA7,L5PHID15_L6PHID30,L2PHIJ7_L3PHIJ7,L5PHID13_L6PHID25,L2PHIK9_L3PHIK9,L1PHIC12_L2PHIB13,L1PHID14_L2PHIB12,L1PHIG25_L2PHIC24,L5PHIB7_L6PHIB10,L3PHID14_L4PHID28,L1PHIF23_L2PHIC21,L5PHID13_L6PHIC22,L2PHIK9_L3PHIK10,L5PHIA4_L6PHIB11,L1PHIG27_L2PHID27,L1PHID14_L2PHIB13,L5PHIA4_L6PHIB9,L3PHID13_L4PHIC24,L5PHIB5_L6PHIB9,L5PHIA1_L6PHIA4,L1PHIB7_L2PHIA5,L5PHIA2_L6PHIA2,L5PHIC9_L6PHIC19,L1PHIH30_L2PHID31,L1PHIG28_L2PHID28,L5PHID13_L6PHID28,L1PHIG26_L2PHID25,L5PHIB5_L6PHIA7,L1PHIE19_L2PHIC21,L3PHIB7_L4PHIB14,L2PHIK10_L3PHIK9,L3PHID16_L4PHID31,L5PHIA3_L6PHIA2,L3PHIA3_L4PHIA6,L1PHIH30_L2PHID28,L3PHIB7_L4PHIB12,L5PHIA1_L6PHIA1,L5PHIA3_L6PHIA4,L1PHIC9_L2PHIB10,L3PHID13_L4PHID28,L1PHIH32_L2PHID31,L5PHIB7_L6PHIC17,L1PHIA3_L2PHIA1,L2PHII2_L3PHII1,L1PHIC12_L2PHIB10,L2PHIJ7_L3PHIJ6,L1PHIE17_L2PHIC18,L3PHID15_L4PHID29,L2PHIK10_L3PHIK11,L5PHIA2_L6PHIA7,L1PHIB5_L2PHIA3,L1PHIH30_L2PHID32,L3PHIC12_L4PHID26,L3PHIB6_L4PHIB11,L2PHIL13_L3PHIL14,L1PHIE19_L2PHIC18,L1PHIB6_L2PHIA6,L3PHIC10_L4PHIC19,L1PHIA2_L2PHIA1,L1PHIG26_L2PHIC24,L2PHIJ5_L3PHII4,L3PHID15_L4PHID31,L5PHIB7_L6PHIB11,L2PHIK11_L3PHIK12,L3PHIB8_L4PHIB13,L5PHIB7_L6PHIB13,L5PHIC10_L6PHIC22,L3PHIB6_L4PHIB9,L3PHID16_L4PHID32,L5PHIC10_L6PHIB16,L3PHIA2_L4PHIA3,L2PHIJ8_L3PHIK9,L1PHIC9_L2PHIA8,L5PHIC10_L6PHIC17,L3PHIC9_L4PHIC20,L3PHIB7_L4PHIB13,L5PHIB7_L6PHIB12,L5PHIA3_L6PHIB9,L5PHIA3_L6PHIA7,L1PHIH31_L2PHID32,L5PHIC9_L6PHIB16,L1PHIA3_L2PHIA5,L1PHIF24_L2PHID25,L3PHID16_L4PHID29,L3PHIB8_L4PHIC18,L1PHID15_L2PHIB15,L3PHIB5_L4PHIB11,L1PHIH31_L2PHID31,L5PHIA4_L6PHIB10,L3PHIC11_L4PHIC23,L3PHIA2_L4PHIA6,L1PHID14_L2PHIB15,L1PHID13_L2PHIB11,L3PHIB7_L4PHIB16,L1PHIE19_L2PHIC19,L5PHIB5_L6PHIA6,L3PHID14_L4PHID26,L1PHIB7_L2PHIA8,L1PHIC10_L2PHIB12,L3PHIC10_L4PHIC17,L1PHIG26_L2PHID26,L5PHIC9_L6PHIC20,L5PHIC9_L6PHIB14,L5PHID16_L6PHID30,L1PHIB8_L2PHIB9,L1PHIE20_L2PHIC18,L3PHIA3_L4PHIA8,L3PHIC11_L4PHIC22,L1PHIH29_L2PHID31,L3PHIB8_L4PHIC17,L1PHIA4_L2PHIA2,L3PHID15_L4PHID28,L1PHIF22_L2PHIC20,L1PHIE17_L2PHIC19,L5PHIB6_L6PHIB14,L1PHIF22_L2PHIC22,L2PHIJ6_L3PHIJ7,L1PHIH30_L2PHID29,L5PHIA2_L6PHIA6,L5PHIB5_L6PHIB13,L5PHIA4_L6PHIA7,L5PHIB5_L6PHIB11,L2PHIL16_L3PHIL16,L5PHIC11_L6PHIC21,L3PHIA4_L4PHIB9,L5PHID14_L6PHID25,L5PHIC10_L6PHIC19,L5PHID14_L6PHID29,L2PHIL16_L3PHIL15,L1PHIC11_L2PHIB10,L1PHID15_L2PHIB16,L1PHIG27_L2PHID25,L3PHIB5_L4PHIB9,L3PHID13_L4PHID27,L3PHIB6_L4PHIB14,L5PHID14_L6PHID27,L3PHIC11_L4PHIC19,L5PHIC12_L6PHID26,L1PHIE20_L2PHIC21,L1PHIB8_L2PHIA8,L2PHIJ8_L3PHIJ7,L1PHIF21_L2PHIC19,L2PHIK9_L3PHIJ8,L2PHIL13_L3PHIK12,L3PHIC9_L4PHIB16,L5PHIC11_L6PHIC22,L3PHIA1_L4PHIA2,L1PHIA3_L2PHIA3,L2PHIL14_L3PHIL13,L3PHIB5_L4PHIB10,L3PHID15_L4PHID30,L1PHIB5_L2PHIA5,L1PHID16_L2PHIC18,L1PHIH31_L2PHID30,L1PHIA2_L2PHIA4,L5PHID15_L6PHID32,L3PHID14_L4PHID27,L2PHIJ7_L3PHIJ8,L5PHIA1_L6PHIA3,L1PHIC10_L2PHIA8,L1PHIB6_L2PHIA7,L5PHIA2_L6PHIA1,L5PHIA4_L6PHIA5,L1PHIF24_L2PHID26,L2PHII1_L3PHII1,L5PHIA2_L6PHIA3,L5PHIB5_L6PHIB10,L3PHIA4_L4PHIB10,L3PHIC10_L4PHIC22,L3PHIA2_L4PHIA4,L2PHIL15_L3PHIL15,L1PHIF21_L2PHIC20,L1PHIA1_L2PHIA1,L3PHIB7_L4PHIB15,L1PHIE17_L2PHIC17,L5PHIB6_L6PHIA8,L1PHIF22_L2PHIC21,L1PHIE20_L2PHIC22,L5PHIC9_L6PHIB15,L1PHIG27_L2PHID26,L5PHIC10_L6PHIC21,L1PHIG28_L2PHID26,L2PHIJ8_L3PHIJ8,L5PHIC11_L6PHIC19,L1PHIC10_L2PHIB10,L2PHIJ6_L3PHIJ5,L1PHIG25_L2PHIC23,L1PHID16_L2PHIB16,L3PHIB6_L4PHIB12,L3PHIB8_L4PHIB15,L1PHIC11_L2PHIB9,L3PHIC9_L4PHIB15,L1PHIE20_L2PHIC20,L1PHIB6_L2PHIA5,L1PHIC11_L2PHIB13,L1PHIC11_L2PHIB11,L5PHIB5_L6PHIA8,L2PHIL15_L3PHIL16,L3PHID14_L4PHID30,L1PHIB6_L2PHIA8,L1PHID16_L2PHIC17,L1PHID15_L2PHIB13,L1PHIF22_L2PHIC24,L1PHIB7_L2PHIA6,L3PHID15_L4PHID27,L1PHIH29_L2PHID27,L5PHIB8_L6PHIB15,L3PHIB5_L4PHIB12,L2PHIJ6_L3PHIJ6,L5PHIA1_L6PHIA5,L1PHIE20_L2PHIC19,L3PHIC12_L4PHID25,L5PHIB6_L6PHIB15,L1PHID13_L2PHIB14,L5PHIB7_L6PHIB15,L2PHIL14_L3PHIL14,L5PHIC11_L6PHIC24,L2PHII2_L3PHII3,L1PHIB8_L2PHIA7,L1PHID13_L2PHIB15,L5PHIC9_L6PHIC17,L5PHID15_L6PHID26,L5PHIA2_L6PHIA4,L3PHIB8_L4PHIB16,L2PHIL13_L3PHIL13,L1PHIA2_L2PHIA3,L3PHIC12_L4PHIC24,L5PHIB6_L6PHIB11,L1PHIB5_L2PHIA4,L5PHIA3_L6PHIA8,L5PHIB7_L6PHIB14,L2PHIK12_L3PHIK11,L1PHIH29_L2PHID30,L3PHID13_L4PHIC23,L1PHIC12_L2PHIB14,L5PHID14_L6PHID30,L1PHIH29_L2PHID29,L1PHIF23_L2PHIC22,L5PHID16_L6PHID31,L2PHII4_L3PHIJ5,L5PHIA3_L6PHIA3,L3PHIB6_L4PHIB13,L1PHID14_L2PHIB16,L5PHIC9_L6PHIC18,L1PHIB6_L2PHIA4,L5PHIC12_L6PHID25,L5PHIB7_L6PHIB16,L1PHIA4_L2PHIA3,L3PHIA2_L4PHIA5,L5PHIA2_L6PHIA5,L2PHIJ5_L3PHIJ6);

  type enum_TPROJ_60 is (L5L6C_L1PHIC,L2L3C_L1PHIE,L5L6A_L2PHIA,L5L6A_L1PHIA,L3L4C_L2PHIC,L5L6B_L2PHIB,L3L4B_L1PHIE,L3L4D_L2PHID,L3L4C_L1PHIG,L1L2K_L3PHID,L3L4B_L1PHID,L5L6C_L1PHIF,L5L6C_L1PHIE,L3L4B_L2PHIA,L2L3C_L1PHIF,L1L2J_L3PHID,L5L6B_L1PHID,L1L2J_L3PHIC,L1L2I_L3PHID,L1L2E_L3PHIB,L2L3A_L1PHIC,L5L6B_L1PHIF,L5L6A_L1PHID,L3L4C_L1PHIE,L5L6C_L2PHID,L1L2G_L3PHIC,L3L4B_L2PHIC,L3L4B_L1PHIC,L2L3D_L1PHIH,L5L6B_L1PHIC,L1L2F_L3PHIB,L1L2D_L3PHIA,L3L4D_L2PHIC,L3L4A_L1PHIB,L1L2F_L3PHIC,L1L2I_L3PHIC,L2L3D_L1PHIG,L3L4A_L1PHIC,L3L4A_L2PHIB,L1L2H_L3PHIC,L5L6A_L1PHIC,L5L6A_L3PHIA,L5L6D_L2PHID,L5L6D_L1PHIE,L5L6D_L1PHIH,L5L6B_L1PHIB,L1L2C_L3PHIA,L5L6B_L2PHIC,L3L4B_L1PHIB,L2L3A_L1PHIB,L2L3B_L1PHIC,L5L6B_L3PHIA,L2L3B_L1PHIE,L3L4D_L1PHIH,L1L2A_L3PHIA,L2L3C_L1PHID,L3L4A_L1PHIA,L5L6D_L1PHIF,L2L3C_L1PHIG,L1L2B_L3PHIB,L5L6B_L3PHIC,L2L3A_L1PHIA,L5L6D_L3PHIC,L5L6B_L2PHIA,L1L2G_L3PHIB,L3L4B_L2PHIB,L1L2L_L3PHID,L5L6B_L3PHIB,L5L6A_L3PHIB,L5L6A_L1PHIB,L5L6C_L3PHIB,L5L6D_L3PHID,L2L3D_L1PHIF,L5L6C_L3PHID,L5L6B_L1PHIE,L5L6C_L3PHIC,L1L2B_L3PHIA,L5L6C_L1PHID,L3L4C_L1PHIF,L1L2D_L3PHIB,L1L2C_L3PHIB,L3L4C_L2PHIB,L5L6C_L2PHIC,L3L4C_L2PHID,L2L3B_L1PHID,L5L6C_L2PHIB,L3L4A_L2PHIA,L3L4D_L1PHIG,L5L6D_L2PHIC,L5L6C_L1PHIG,L5L6D_L1PHIG,L3L4C_L1PHID,L5L6A_L2PHIB,L3L4D_L1PHIF);

  type enum_TPROJ_58 is (L2L3C_L5PHIB,L1L2E_L5PHIC,L1L2H_L6PHIC,L3L4B_L5PHIA,L3L4C_L5PHIB,L1L2L_L6PHIC,L1L2H_L4PHIB,L1L2H_L5PHID,L1L2L_L4PHID,L2L3C_L5PHID,L1L2H_L6PHID,L1L2E_L6PHIB,L1L2J_L6PHID,L1L2L_L5PHID,L1L2K_L4PHID,L1L2H_L4PHIC,L3L4B_L5PHIC,L1L2K_L4PHIC,L1L2G_L4PHIC,L3L4D_L6PHIC,L5L6A_L4PHIA,L3L4C_L5PHID,L1L2A_L5PHIB,L2L3B_L5PHIB,L1L2C_L6PHIB,L3L4D_L6PHID,L5L6A_L4PHIB,L5L6D_L4PHID,L1L2G_L6PHID,L2L3D_L4PHID,L1L2D_L5PHIC,L1L2I_L5PHID,L1L2E_L4PHIC,L1L2E_L4PHIA,L2L3B_L4PHIA,L1L2I_L4PHIC,L1L2I_L4PHID,L1L2G_L6PHIB,L2L3D_L5PHIC,L1L2F_L5PHIC,L2L3A_L4PHIA,L5L6C_L4PHIB,L1L2B_L5PHIA,L1L2G_L4PHIB,L1L2F_L6PHIA,L1L2H_L5PHIB,L2L3B_L5PHIC,L1L2H_L5PHIC,L1L2J_L5PHID,L1L2D_L4PHIA,L1L2D_L6PHIB,L1L2I_L5PHIB,L1L2A_L4PHIA,L1L2D_L6PHIA,L1L2C_L4PHIA,L3L4A_L6PHIA,L1L2A_L6PHIB,L2L3A_L5PHIA,L3L4D_L5PHID,L1L2E_L4PHIB,L5L6B_L4PHIC,L2L3D_L5PHID,L1L2C_L5PHIA,L1L2I_L6PHID,L3L4C_L6PHIB,L3L4C_L6PHIC,L2L3A_L5PHIB,L1L2J_L5PHIC,L1L2B_L4PHIA,L3L4A_L5PHIA,L1L2A_L5PHIA,L3L4B_L6PHIA,L1L2C_L4PHIB,L1L2B_L6PHIB,L1L2B_L4PHIB,L2L3D_L4PHIC,L1L2G_L5PHIC,L1L2E_L6PHIA,L5L6B_L4PHIB,L1L2G_L6PHIC,L3L4B_L5PHIB,L2L3A_L4PHIB,L1L2I_L6PHIC,L1L2C_L6PHIA,L2L3B_L4PHIB,L1L2J_L4PHID,L1L2F_L5PHIB,L1L2D_L6PHIC,L1L2K_L6PHIC,L1L2H_L6PHIB,L1L2K_L5PHIC,L3L4C_L6PHID,L1L2K_L6PHID,L2L3C_L4PHIB,L1L2L_L5PHIC,L5L6C_L4PHIC,L3L4A_L6PHIB,L1L2D_L5PHIA,L1L2F_L4PHIC,L1L2J_L4PHIC,L1L2J_L6PHIC,L1L2E_L5PHIA,L1L2B_L5PHIB,L1L2I_L6PHIB,L2L3C_L4PHIC,L1L2E_L5PHIB,L1L2G_L5PHIB,L3L4C_L5PHIC,L3L4A_L5PHIB,L1L2E_L6PHIC,L1L2C_L5PHIB,L5L6B_L4PHIA,L2L3B_L5PHIA,L2L3C_L4PHID,L1L2B_L6PHIA,L1L2I_L5PHIC,L5L6D_L4PHIC,L2L3C_L5PHIC,L1L2H_L4PHID,L1L2F_L6PHIC,L1L2F_L6PHIB,L3L4B_L6PHIC,L5L6C_L4PHID,L1L2D_L5PHIB,L1L2F_L4PHIB,L1L2K_L5PHID,L1L2D_L4PHIB,L2L3B_L4PHIC,L3L4B_L6PHIB,L3L4D_L5PHIC);

  type enum_TPAR_70 is (L1L2F,L1L2I,L1L2D,L2L3B,L3L4D,L3L4A,L3L4C,L5L6C,L1L2E,L5L6A,L2L3D,L1L2C,L1L2J,L5L6B,L1L2B,L2L3A,L1L2K,L1L2L,L1L2H,L2L3C,L1L2G,L3L4B,L5L6D,L1L2A);

  type enum_VMPROJ_24 is (L4PHIB16,L2PHID26,L4PHID32,L4PHID25,L5PHIC22,L3PHIC24,L4PHIA5,L6PHID28,L6PHIB11,L2PHIB10,L1PHIA4,L3PHIC17,L2PHID25,L6PHID26,L1PHIC10,L2PHID28,L6PHID31,L6PHIA3,L2PHIC19,L1PHID16,L3PHID26,L3PHID28,L4PHIA7,L4PHIC19,L1PHID14,L3PHIC21,L6PHIA2,L5PHIA7,L6PHIB13,L4PHIA3,L4PHIA4,L4PHIC24,L5PHIB9,L3PHIA5,L4PHIB12,L3PHIC18,L5PHIA5,L1PHIE19,L3PHIC19,L3PHIA8,L2PHIA7,L6PHIB15,L5PHIB12,L4PHIC20,L2PHIB14,L1PHIG28,L1PHIB5,L3PHIB11,L6PHIC23,L5PHID32,L2PHIA5,L3PHIB16,L2PHIB15,L5PHIA8,L2PHIA3,L1PHIH31,L1PHIC11,L1PHIB6,L2PHIB9,L1PHIH32,L1PHIG27,L4PHIB9,L2PHIA8,L5PHID27,L6PHIA8,L3PHID25,L5PHIB15,L1PHIH29,L4PHID30,L3PHIC22,L6PHID29,L5PHIA4,L1PHID15,L5PHID30,L4PHID31,L6PHIC20,L6PHIA4,L4PHID26,L5PHIC21,L2PHIC23,L4PHIA8,L5PHID29,L3PHID29,L4PHIB14,L4PHIA6,L3PHIB10,L2PHIA1,L4PHIB11,L5PHIA2,L6PHIC17,L1PHIA2,L3PHID27,L1PHIF21,L6PHIB9,L5PHIC17,L5PHIA6,L1PHIF23,L5PHID28,L1PHIB8,L3PHIA1,L5PHID26,L5PHIC20,L1PHID13,L2PHIC18,L3PHIA7,L6PHIC18,L6PHIC21,L4PHIC22,L2PHID32,L3PHID32,L6PHID27,L1PHIC9,L5PHIA3,L2PHIB13,L2PHIC17,L4PHIB15,L1PHIA1,L6PHIA5,L5PHIB10,L1PHIC12,L4PHIA1,L1PHIE17,L3PHID31,L2PHIA6,L3PHIA4,L2PHIC20,L6PHIB16,L1PHIB7,L2PHID29,L6PHID32,L4PHIC21,L4PHIB10,L3PHIA6,L6PHID30,L3PHIB12,L5PHIB14,L5PHIC23,L5PHIC24,L6PHIB10,L2PHIC24,L4PHID28,L5PHIA1,L6PHIC22,L4PHIC17,L3PHIB14,L5PHID25,L2PHIA4,L5PHIC19,L6PHIC24,L6PHIB12,L4PHIB13,L6PHIA1,L6PHIA6,L2PHID31,L3PHIB15,L4PHID27,L1PHIA3,L2PHIC22,L6PHIC19,L2PHIA2,L1PHIG25,L4PHIC23,L2PHIC21,L6PHIB14,L6PHID25,L1PHIF22,L2PHID27,L4PHIC18,L1PHIF24,L3PHIB13,L1PHIH30,L3PHIC20,L2PHIB16,L2PHIB12,L3PHID30,L1PHIE18,L5PHIC18,L2PHID30,L6PHIA7,L5PHIB11,L3PHIA3,L1PHIE20,L5PHIB16,L5PHID31,L4PHID29,L4PHIA2,L5PHIB13,L1PHIG26,L3PHIB9,L2PHIB11,L3PHIC23,L3PHIA2);

  type enum_AP_60 is (L1PHIG,L1PHIA,L2PHID,L3PHIB,L2PHIC,L3PHIC,L3PHIA,L1PHIH,L1PHIE,L1PHIF,L1PHID,L3PHID,L1PHIB,L2PHIB,L1PHIC,L2PHIA);

  type enum_AP_58 is (L4PHIA,L5PHIA,L5PHIB,L6PHIC,L6PHIB,L4PHIC,L4PHID,L4PHIB,L6PHID,L5PHIC,L6PHIA,L5PHID);

  type enum_CM_14 is (L5PHIC17,L5PHIA5,L4PHID28,L1PHID15,L1PHIB6,L2PHID26,L4PHID25,L2PHIB15,L3PHIC20,L1PHIF22,L2PHIA4,L1PHIA1,L3PHIC23,L2PHID25,L2PHID27,L5PHIB13,L3PHIB9,L6PHIC18,L4PHIB11,L6PHIB15,L1PHIH29,L2PHID31,L1PHID16,L3PHID26,L5PHIC24,L1PHIE17,L1PHIB7,L2PHID29,L3PHIA4,L3PHIC22,L4PHIB14,L3PHID28,L2PHIC23,L5PHID29,L3PHIB12,L6PHIB13,L2PHIC21,L5PHIA6,L2PHIC19,L4PHIB12,L1PHIB5,L3PHIC24,L5PHIA7,L2PHIA3,L4PHID31,L2PHIB12,L1PHIE18,L3PHIB11,L6PHIC20,L5PHIC20,L5PHID25,L6PHIB11,L4PHIC17,L4PHIC21,L1PHIC11,L3PHIA2,L1PHID14,L5PHIB14,L6PHID30,L3PHIC18,L3PHID25,L2PHID32,L4PHIA7,L1PHIF21,L6PHIB10,L6PHIB9,L4PHIC22,L2PHIB10,L1PHID13,L5PHIA2,L6PHIA7,L3PHIC21,L1PHIC12,L6PHID25,L5PHIB16,L5PHID32,L6PHID27,L6PHIB12,L4PHIA6,L2PHIC22,L5PHIC19,L2PHIC18,L6PHIC24,L2PHIA2,L4PHIC19,L5PHIA3,L2PHIB13,L6PHIA8,L6PHID32,L6PHIA2,L5PHIA4,L3PHIA8,L5PHIC21,L5PHIC18,L5PHIB9,L1PHIG26,L5PHIA1,L5PHID30,L6PHIC23,L5PHIB10,L4PHIA5,L3PHIB14,L4PHID30,L6PHIC19,L2PHIA1,L3PHIA6,L1PHIF24,L4PHIB10,L4PHIA8,L3PHID30,L5PHIB12,L3PHID27,L3PHIB10,L4PHIC20,L5PHID27,L4PHID29,L1PHIH30,L4PHIB16,L1PHIG28,L3PHIB13,L1PHIC9,L6PHIA1,L4PHID27,L1PHIA4,L6PHID28,L2PHIC24,L2PHIA7,L4PHIA4,L4PHIB15,L2PHIB14,L4PHIB13,L1PHIH31,L3PHIA7,L6PHID31,L3PHIA1,L6PHID26,L5PHIC22,L6PHIC21,L2PHIC17,L5PHID28,L4PHIC24,L2PHIA6,L5PHIB11,L3PHIB16,L2PHIA8,L5PHID26,L4PHID32,L2PHIA5,L4PHID26,L1PHIC10,L2PHID28,L1PHIE20,L2PHID30,L4PHIC18,L2PHIC20,L6PHIB14,L3PHID32,L3PHIB15,L4PHIB9,L1PHIB8,L2PHIB9,L6PHIC22,L5PHIB15,L3PHIA3,L3PHID29,L6PHIC17,L1PHIH32,L1PHIE19,L4PHIA3,L5PHID31,L3PHIA5,L4PHIA1,L6PHID29,L1PHIA2,L5PHIC23,L1PHIA3,L6PHIA4,L4PHIC23,L2PHIB16,L1PHIG25,L2PHIB11,L6PHIA3,L3PHIC19,L3PHID31,L4PHIA2,L6PHIA5,L5PHIA8,L6PHIA6,L1PHIG27,L1PHIF23,L3PHIC17,L6PHIB16);

  type enum_FM_52 is (L5L6_L1PHIF,L2L3_L1PHIG,L2L3_L1PHID,L3L4_L5PHIB,L3L4_L1PHIA,L3L4_L1PHIC,L1L2_L6PHIA,L2L3_L5PHIB,L2L3_L5PHIA,L1L2_L3PHIA,L3L4_L2PHID,L1L2_L5PHIC,L2L3_L4PHIA,L3L4_L1PHIH,L5L6_L2PHIA,L5L6_L3PHID,L3L4_L1PHIB,L5L6_L4PHID,L1L2_L5PHIA,L1L2_L4PHID,L2L3_L5PHID,L5L6_L2PHIB,L1L2_L3PHID,L2L3_L4PHIB,L1L2_L3PHIB,L5L6_L3PHIA,L2L3_L1PHIC,L3L4_L1PHIF,L3L4_L2PHIA,L3L4_L6PHIB,L2L3_L4PHID,L1L2_L4PHIB,L3L4_L1PHID,L5L6_L1PHID,L3L4_L1PHIG,L3L4_L1PHIE,L2L3_L1PHIB,L1L2_L3PHIC,L2L3_L1PHIH,L5L6_L4PHIC,L3L4_L2PHIB,L5L6_L1PHIG,L1L2_L4PHIC,L3L4_L2PHIC,L2L3_L1PHIF,L1L2_L4PHIA,L3L4_L5PHIA,L1L2_L5PHIB,L5L6_L4PHIA,L1L2_L6PHIC,L3L4_L5PHID,L2L3_L1PHIA,L1L2_L5PHID,L3L4_L6PHID,L5L6_L1PHIA,L5L6_L3PHIC,L1L2_L6PHIB,L5L6_L1PHIH,L5L6_L1PHIC,L5L6_L1PHIB,L3L4_L6PHIA,L5L6_L1PHIE,L3L4_L6PHIC,L2L3_L1PHIE,L5L6_L4PHIB,L2L3_L4PHIC,L3L4_L5PHIC,L2L3_L5PHIC,L5L6_L2PHID,L1L2_L6PHID,L5L6_L2PHIC,L5L6_L3PHIB);

  type enum_TW_84 is (L5L6,L1L2,L3L4,L2L3);

  type enum_BW_46 is (L5L6_L1,L5L6_L2,L5L6_L3,L5L6_L4,L1L2_L3,L1L2_L4,L1L2_L5,L1L2_L6,L3L4_L1,L3L4_L2,L3L4_L5,L3L4_L6,L2L3_L1,L2L3_L4,L2L3_L5);

  type t_arr_DL_39_1b is array(enum_DL_39) of std_logic;
  type t_arr_DL_39_DATA is array(enum_DL_39) of std_logic_vector(38 downto 0);
  type t_arr_IL_36_1b is array(enum_IL_36) of std_logic;
  type t_arr_IL_36_ADDR is array(enum_IL_36) of std_logic_vector(7 downto 0);
  type t_arr_IL_36_DATA is array(enum_IL_36) of std_logic_vector(35 downto 0);
  type t_arr_IL_36_NENT is array(enum_IL_36) of t_arr2_7b;
  type t_arr_AS_36_1b is array(enum_AS_36) of std_logic;
  type t_arr_AS_36_ADDR is array(enum_AS_36) of std_logic_vector(9 downto 0);
  type t_arr_AS_36_DATA is array(enum_AS_36) of std_logic_vector(35 downto 0);
  type t_arr_AS_36_NENT is array(enum_AS_36) of t_arr8_7b;
  type t_arr_VMSME_17_1b is array(enum_VMSME_17) of std_logic;
  type t_arr_VMSME_17_ADDR is array(enum_VMSME_17) of std_logic_vector(9 downto 0);
  type t_arr_VMSME_17_DATA is array(enum_VMSME_17) of std_logic_vector(16 downto 0);
  type t_arr_VMSME_17_NENT is array(enum_VMSME_17) of t_arr8_8_5b;
  type t_arr_VMSME_16_1b is array(enum_VMSME_16) of std_logic;
  type t_arr_VMSME_16_ADDR is array(enum_VMSME_16) of std_logic_vector(9 downto 0);
  type t_arr_VMSME_16_DATA is array(enum_VMSME_16) of std_logic_vector(15 downto 0);
  type t_arr_VMSME_16_NENT is array(enum_VMSME_16) of t_arr8_8_5b;
  type t_arr_VMSTE_22_1b is array(enum_VMSTE_22) of std_logic;
  type t_arr_VMSTE_22_ADDR is array(enum_VMSTE_22) of std_logic_vector(7 downto 0);
  type t_arr_VMSTE_22_DATA is array(enum_VMSTE_22) of std_logic_vector(21 downto 0);
  type t_arr_VMSTE_22_NENT is array(enum_VMSTE_22) of t_arr2_7b;
  type t_arr_VMSTE_17_1b is array(enum_VMSTE_17) of std_logic;
  type t_arr_VMSTE_17_ADDR is array(enum_VMSTE_17) of std_logic_vector(7 downto 0);
  type t_arr_VMSTE_17_DATA is array(enum_VMSTE_17) of std_logic_vector(16 downto 0);
  type t_arr_VMSTE_17_NENT is array(enum_VMSTE_17) of t_arr2_8_5b;
  type t_arr_VMSTE_23_1b is array(enum_VMSTE_23) of std_logic;
  type t_arr_VMSTE_23_ADDR is array(enum_VMSTE_23) of std_logic_vector(7 downto 0);
  type t_arr_VMSTE_23_DATA is array(enum_VMSTE_23) of std_logic_vector(22 downto 0);
  type t_arr_VMSTE_23_NENT is array(enum_VMSTE_23) of t_arr2_7b;
  type t_arr_VMSTE_16_1b is array(enum_VMSTE_16) of std_logic;
  type t_arr_VMSTE_16_ADDR is array(enum_VMSTE_16) of std_logic_vector(7 downto 0);
  type t_arr_VMSTE_16_DATA is array(enum_VMSTE_16) of std_logic_vector(15 downto 0);
  type t_arr_VMSTE_16_NENT is array(enum_VMSTE_16) of t_arr2_8_5b;
  type t_arr_SP_14_1b is array(enum_SP_14) of std_logic;
  type t_arr_SP_14_ADDR is array(enum_SP_14) of std_logic_vector(7 downto 0);
  type t_arr_SP_14_DATA is array(enum_SP_14) of std_logic_vector(13 downto 0);
  type t_arr_SP_14_NENT is array(enum_SP_14) of t_arr2_7b;
  type t_arr_TPROJ_60_1b is array(enum_TPROJ_60) of std_logic;
  type t_arr_TPROJ_60_ADDR is array(enum_TPROJ_60) of std_logic_vector(7 downto 0);
  type t_arr_TPROJ_60_DATA is array(enum_TPROJ_60) of std_logic_vector(59 downto 0);
  type t_arr_TPROJ_60_NENT is array(enum_TPROJ_60) of t_arr2_7b;
  type t_arr_TPROJ_58_1b is array(enum_TPROJ_58) of std_logic;
  type t_arr_TPROJ_58_ADDR is array(enum_TPROJ_58) of std_logic_vector(7 downto 0);
  type t_arr_TPROJ_58_DATA is array(enum_TPROJ_58) of std_logic_vector(57 downto 0);
  type t_arr_TPROJ_58_NENT is array(enum_TPROJ_58) of t_arr2_7b;
  type t_arr_TPAR_70_1b is array(enum_TPAR_70) of std_logic;
  type t_arr_TPAR_70_ADDR is array(enum_TPAR_70) of std_logic_vector(9 downto 0);
  type t_arr_TPAR_70_DATA is array(enum_TPAR_70) of std_logic_vector(69 downto 0);
  type t_arr_TPAR_70_NENT is array(enum_TPAR_70) of t_arr8_7b;
  type t_arr_VMPROJ_24_1b is array(enum_VMPROJ_24) of std_logic;
  type t_arr_VMPROJ_24_ADDR is array(enum_VMPROJ_24) of std_logic_vector(7 downto 0);
  type t_arr_VMPROJ_24_DATA is array(enum_VMPROJ_24) of std_logic_vector(23 downto 0);
  type t_arr_VMPROJ_24_NENT is array(enum_VMPROJ_24) of t_arr2_7b;
  type t_arr_AP_60_1b is array(enum_AP_60) of std_logic;
  type t_arr_AP_60_ADDR is array(enum_AP_60) of std_logic_vector(9 downto 0);
  type t_arr_AP_60_DATA is array(enum_AP_60) of std_logic_vector(59 downto 0);
  type t_arr_AP_60_NENT is array(enum_AP_60) of t_arr8_7b;
  type t_arr_AP_58_1b is array(enum_AP_58) of std_logic;
  type t_arr_AP_58_ADDR is array(enum_AP_58) of std_logic_vector(9 downto 0);
  type t_arr_AP_58_DATA is array(enum_AP_58) of std_logic_vector(57 downto 0);
  type t_arr_AP_58_NENT is array(enum_AP_58) of t_arr8_7b;
  type t_arr_CM_14_1b is array(enum_CM_14) of std_logic;
  type t_arr_CM_14_ADDR is array(enum_CM_14) of std_logic_vector(7 downto 0);
  type t_arr_CM_14_DATA is array(enum_CM_14) of std_logic_vector(13 downto 0);
  type t_arr_CM_14_NENT is array(enum_CM_14) of t_arr2_7b;
  type t_arr_FM_52_1b is array(enum_FM_52) of std_logic;
  type t_arr_FM_52_ADDR is array(enum_FM_52) of std_logic_vector(7 downto 0);
  type t_arr_FM_52_DATA is array(enum_FM_52) of std_logic_vector(51 downto 0);
  type t_arr_FM_52_NENT is array(enum_FM_52) of t_arr2_7b;
  type t_arr_TW_84_1b is array(enum_TW_84) of std_logic;
  type t_arr_TW_84_DATA is array(enum_TW_84) of std_logic_vector(83 downto 0);
  type t_arr_BW_46_1b is array(enum_BW_46) of std_logic;
  type t_arr_BW_46_DATA is array(enum_BW_46) of std_logic_vector(45 downto 0);

  -- ########################### Functions ###########################

  -- Following functions are needed because VHDL doesn't preserve case when converting an enum to a string using image
  function memory_enum_to_string(val: enum_DL_39) return string;
  function memory_enum_to_string(val: enum_IL_36) return string;
  function memory_enum_to_string(val: enum_AS_36) return string;
  function memory_enum_to_string(val: enum_VMSME_17) return string;
  function memory_enum_to_string(val: enum_VMSME_16) return string;
  function memory_enum_to_string(val: enum_VMSTE_22) return string;
  function memory_enum_to_string(val: enum_VMSTE_17) return string;
  function memory_enum_to_string(val: enum_VMSTE_23) return string;
  function memory_enum_to_string(val: enum_VMSTE_16) return string;
  function memory_enum_to_string(val: enum_SP_14) return string;
  function memory_enum_to_string(val: enum_TPROJ_60) return string;
  function memory_enum_to_string(val: enum_TPROJ_58) return string;
  function memory_enum_to_string(val: enum_TPAR_70) return string;
  function memory_enum_to_string(val: enum_VMPROJ_24) return string;
  function memory_enum_to_string(val: enum_AP_60) return string;
  function memory_enum_to_string(val: enum_AP_58) return string;
  function memory_enum_to_string(val: enum_CM_14) return string;
  function memory_enum_to_string(val: enum_FM_52) return string;
  function memory_enum_to_string(val: enum_TW_84) return string;
  function memory_enum_to_string(val: enum_BW_46) return string;

end package memUtil_pkg;

package body memUtil_pkg is

  -- ########################### Functions ###########################

  function memory_enum_to_string(val: enum_DL_39) return string is
  begin
    case val is
       when negPS10G_2_A => return "negPS10G_2_A";
       when neg2S_3_A => return "neg2S_3_A";
       when negPS_1_A => return "negPS_1_A";
       when PS10G_2_A => return "PS10G_2_A";
       when neg2S_4_B => return "neg2S_4_B";
       when negPS_2_A => return "negPS_2_A";
       when twoS_2_B => return "2S_2_B";
       when twoS_4_B => return "2S_4_B";
       when PS10G_3_A => return "PS10G_3_A";
       when twoS_2_A => return "2S_2_A";
       when PS10G_1_A => return "PS10G_1_A";
       when PS_1_A => return "PS_1_A";
       when neg2S_4_A => return "neg2S_4_A";
       when twoS_1_B => return "2S_1_B";
       when negPS10G_1_A => return "negPS10G_1_A";
       when PS_1_B => return "PS_1_B";
       when twoS_3_B => return "2S_3_B";
       when PS10G_2_B => return "PS10G_2_B";
       when negPS10G_3_A => return "negPS10G_3_A";
       when PS10G_1_B => return "PS10G_1_B";
       when neg2S_1_B => return "neg2S_1_B";
       when neg2S_1_A => return "neg2S_1_A";
       when negPS_1_B => return "negPS_1_B";
       when neg2S_2_B => return "neg2S_2_B";
       when PS10G_3_B => return "PS10G_3_B";
       when PS_2_A => return "PS_2_A";
       when neg2S_3_B => return "neg2S_3_B";
       when twoS_1_A => return "2S_1_A";
       when negPS10G_3_B => return "negPS10G_3_B";
       when negPS10G_2_B => return "negPS10G_2_B";
       when PS_2_B => return "PS_2_B";
       when neg2S_2_A => return "neg2S_2_A";
       when negPS_2_B => return "negPS_2_B";
       when negPS10G_1_B => return "negPS10G_1_B";
       when twoS_3_A => return "2S_3_A";
       when twoS_4_A => return "2S_4_A";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_IL_36) return string is
  begin
    case val is
       when L1PHIH_PS10G_2_B => return "L1PHIH_PS10G_2_B";
       when L3PHIB_negPS_2_B => return "L3PHIB_negPS_2_B";
       when L6PHIB_neg2S_4_A => return "L6PHIB_neg2S_4_A";
       when L1PHID_PS10G_1_A => return "L1PHID_PS10G_1_A";
       when L6PHIC_neg2S_3_B => return "L6PHIC_neg2S_3_B";
       when L6PHIC_neg2S_4_B => return "L6PHIC_neg2S_4_B";
       when L2PHIC_PS10G_3_A => return "L2PHIC_PS10G_3_A";
       when L1PHIH_negPS10G_2_B => return "L1PHIH_negPS10G_2_B";
       when L1PHID_PS10G_2_A => return "L1PHID_PS10G_2_A";
       when L3PHIA_negPS_1_A => return "L3PHIA_negPS_1_A";
       when L5PHID_2S_2_B => return "L5PHID_2S_2_B";
       when L5PHIC_neg2S_1_B => return "L5PHIC_neg2S_1_B";
       when L2PHIB_negPS10G_3_A => return "L2PHIB_negPS10G_3_A";
       when L6PHIB_2S_3_B => return "L6PHIB_2S_3_B";
       when L1PHIF_negPS10G_2_B => return "L1PHIF_negPS10G_2_B";
       when L5PHIC_neg2S_2_B => return "L5PHIC_neg2S_2_B";
       when L4PHIC_neg2S_1_B => return "L4PHIC_neg2S_1_B";
       when L3PHID_PS_2_B => return "L3PHID_PS_2_B";
       when L6PHIC_2S_3_B => return "L6PHIC_2S_3_B";
       when L2PHIB_PS10G_3_A => return "L2PHIB_PS10G_3_A";
       when L3PHIA_PS_1_A => return "L3PHIA_PS_1_A";
       when L6PHIB_neg2S_3_A => return "L6PHIB_neg2S_3_A";
       when L5PHIB_neg2S_2_B => return "L5PHIB_neg2S_2_B";
       when L6PHIB_2S_4_A => return "L6PHIB_2S_4_A";
       when L5PHIC_2S_2_A => return "L5PHIC_2S_2_A";
       when L1PHIF_PS10G_1_B => return "L1PHIF_PS10G_1_B";
       when L2PHIA_PS10G_3_A => return "L2PHIA_PS10G_3_A";
       when L1PHIC_negPS10G_2_B => return "L1PHIC_negPS10G_2_B";
       when L6PHIA_2S_3_A => return "L6PHIA_2S_3_A";
       when L1PHIE_PS10G_2_A => return "L1PHIE_PS10G_2_A";
       when L1PHIA_negPS10G_1_A => return "L1PHIA_negPS10G_1_A";
       when L1PHIB_negPS10G_1_A => return "L1PHIB_negPS10G_1_A";
       when L6PHIB_2S_3_A => return "L6PHIB_2S_3_A";
       when L1PHIF_PS10G_2_A => return "L1PHIF_PS10G_2_A";
       when L3PHIB_PS_1_A => return "L3PHIB_PS_1_A";
       when L1PHIH_negPS10G_1_B => return "L1PHIH_negPS10G_1_B";
       when L1PHIE_PS10G_2_B => return "L1PHIE_PS10G_2_B";
       when L5PHIB_neg2S_2_A => return "L5PHIB_neg2S_2_A";
       when L5PHIB_neg2S_1_A => return "L5PHIB_neg2S_1_A";
       when L4PHIA_2S_1_A => return "L4PHIA_2S_1_A";
       when L6PHIC_2S_3_A => return "L6PHIC_2S_3_A";
       when L1PHIF_PS10G_1_A => return "L1PHIF_PS10G_1_A";
       when L5PHIB_2S_2_A => return "L5PHIB_2S_2_A";
       when L3PHID_PS_1_B => return "L3PHID_PS_1_B";
       when L1PHIG_PS10G_2_B => return "L1PHIG_PS10G_2_B";
       when L3PHIC_negPS_2_A => return "L3PHIC_negPS_2_A";
       when L1PHIA_PS10G_1_A => return "L1PHIA_PS10G_1_A";
       when L1PHIC_negPS10G_1_A => return "L1PHIC_negPS10G_1_A";
       when L2PHIB_PS10G_3_B => return "L2PHIB_PS10G_3_B";
       when L3PHID_negPS_2_B => return "L3PHID_negPS_2_B";
       when L1PHIB_PS10G_2_A => return "L1PHIB_PS10G_2_A";
       when L5PHID_neg2S_1_B => return "L5PHID_neg2S_1_B";
       when L4PHIC_2S_1_B => return "L4PHIC_2S_1_B";
       when L1PHIE_negPS10G_1_B => return "L1PHIE_negPS10G_1_B";
       when L2PHIA_negPS10G_3_A => return "L2PHIA_negPS10G_3_A";
       when L1PHID_negPS10G_2_B => return "L1PHID_negPS10G_2_B";
       when L5PHIC_2S_1_B => return "L5PHIC_2S_1_B";
       when L3PHIB_negPS_1_A => return "L3PHIB_negPS_1_A";
       when L5PHIA_neg2S_1_A => return "L5PHIA_neg2S_1_A";
       when L3PHID_negPS_1_B => return "L3PHID_negPS_1_B";
       when L4PHID_2S_1_B => return "L4PHID_2S_1_B";
       when L1PHIC_negPS10G_1_B => return "L1PHIC_negPS10G_1_B";
       when L1PHID_negPS10G_1_B => return "L1PHID_negPS10G_1_B";
       when L1PHIG_PS10G_1_A => return "L1PHIG_PS10G_1_A";
       when L2PHIB_negPS10G_3_B => return "L2PHIB_negPS10G_3_B";
       when L1PHID_PS10G_2_B => return "L1PHID_PS10G_2_B";
       when L1PHIE_PS10G_1_B => return "L1PHIE_PS10G_1_B";
       when L4PHIB_neg2S_1_B => return "L4PHIB_neg2S_1_B";
       when L1PHIF_negPS10G_2_A => return "L1PHIF_negPS10G_2_A";
       when L5PHID_2S_1_B => return "L5PHID_2S_1_B";
       when L1PHIG_PS10G_1_B => return "L1PHIG_PS10G_1_B";
       when L3PHIB_PS_2_A => return "L3PHIB_PS_2_A";
       when L1PHIC_PS10G_1_A => return "L1PHIC_PS10G_1_A";
       when L3PHIC_PS_2_A => return "L3PHIC_PS_2_A";
       when L1PHIG_negPS10G_2_B => return "L1PHIG_negPS10G_2_B";
       when L1PHIF_negPS10G_1_B => return "L1PHIF_negPS10G_1_B";
       when L6PHIA_2S_4_A => return "L6PHIA_2S_4_A";
       when L5PHIC_2S_2_B => return "L5PHIC_2S_2_B";
       when L2PHID_PS10G_3_B => return "L2PHID_PS10G_3_B";
       when L3PHIB_negPS_2_A => return "L3PHIB_negPS_2_A";
       when L6PHID_2S_4_B => return "L6PHID_2S_4_B";
       when L1PHIE_negPS10G_2_B => return "L1PHIE_negPS10G_2_B";
       when L1PHIB_PS10G_1_A => return "L1PHIB_PS10G_1_A";
       when L4PHID_neg2S_1_B => return "L4PHID_neg2S_1_B";
       when L1PHIC_PS10G_2_B => return "L1PHIC_PS10G_2_B";
       when L1PHIC_negPS10G_2_A => return "L1PHIC_negPS10G_2_A";
       when L5PHIA_neg2S_2_A => return "L5PHIA_neg2S_2_A";
       when L4PHIB_neg2S_1_A => return "L4PHIB_neg2S_1_A";
       when L3PHIB_PS_1_B => return "L3PHIB_PS_1_B";
       when L1PHIB_negPS10G_2_A => return "L1PHIB_negPS10G_2_A";
       when L1PHIH_PS10G_1_B => return "L1PHIH_PS10G_1_B";
       when L4PHIC_2S_1_A => return "L4PHIC_2S_1_A";
       when L6PHIB_neg2S_3_B => return "L6PHIB_neg2S_3_B";
       when L3PHIC_PS_2_B => return "L3PHIC_PS_2_B";
       when L3PHIB_PS_2_B => return "L3PHIB_PS_2_B";
       when L6PHID_neg2S_4_B => return "L6PHID_neg2S_4_B";
       when L3PHIA_PS_2_A => return "L3PHIA_PS_2_A";
       when L5PHIB_2S_1_A => return "L5PHIB_2S_1_A";
       when L1PHIF_PS10G_2_B => return "L1PHIF_PS10G_2_B";
       when L5PHIA_2S_1_A => return "L5PHIA_2S_1_A";
       when L3PHIC_PS_1_B => return "L3PHIC_PS_1_B";
       when L4PHIC_neg2S_1_A => return "L4PHIC_neg2S_1_A";
       when L1PHIA_PS10G_2_A => return "L1PHIA_PS10G_2_A";
       when L6PHIB_neg2S_4_B => return "L6PHIB_neg2S_4_B";
       when L1PHID_negPS10G_2_A => return "L1PHID_negPS10G_2_A";
       when L4PHIB_2S_1_B => return "L4PHIB_2S_1_B";
       when L1PHIA_negPS10G_2_A => return "L1PHIA_negPS10G_2_A";
       when L6PHID_neg2S_3_B => return "L6PHID_neg2S_3_B";
       when L6PHIC_2S_4_B => return "L6PHIC_2S_4_B";
       when L2PHIC_negPS10G_3_A => return "L2PHIC_negPS10G_3_A";
       when L6PHIC_neg2S_3_A => return "L6PHIC_neg2S_3_A";
       when L2PHID_negPS10G_3_B => return "L2PHID_negPS10G_3_B";
       when L3PHIC_negPS_1_B => return "L3PHIC_negPS_1_B";
       when L3PHIB_negPS_1_B => return "L3PHIB_negPS_1_B";
       when L3PHIA_negPS_2_A => return "L3PHIA_negPS_2_A";
       when L5PHID_neg2S_2_B => return "L5PHID_neg2S_2_B";
       when L5PHIB_2S_2_B => return "L5PHIB_2S_2_B";
       when L5PHIC_neg2S_2_A => return "L5PHIC_neg2S_2_A";
       when L1PHIE_negPS10G_2_A => return "L1PHIE_negPS10G_2_A";
       when L6PHIB_2S_4_B => return "L6PHIB_2S_4_B";
       when L4PHIB_2S_1_A => return "L4PHIB_2S_1_A";
       when L3PHIC_negPS_2_B => return "L3PHIC_negPS_2_B";
       when L6PHIC_2S_4_A => return "L6PHIC_2S_4_A";
       when L3PHIC_PS_1_A => return "L3PHIC_PS_1_A";
       when L2PHIC_negPS10G_3_B => return "L2PHIC_negPS10G_3_B";
       when L6PHID_2S_3_B => return "L6PHID_2S_3_B";
       when L4PHIA_neg2S_1_A => return "L4PHIA_neg2S_1_A";
       when L1PHIC_PS10G_2_A => return "L1PHIC_PS10G_2_A";
       when L1PHIG_negPS10G_1_B => return "L1PHIG_negPS10G_1_B";
       when L6PHIA_neg2S_4_A => return "L6PHIA_neg2S_4_A";
       when L1PHIE_PS10G_1_A => return "L1PHIE_PS10G_1_A";
       when L6PHIC_neg2S_4_A => return "L6PHIC_neg2S_4_A";
       when L2PHIC_PS10G_3_B => return "L2PHIC_PS10G_3_B";
       when L5PHIA_2S_2_A => return "L5PHIA_2S_2_A";
       when L1PHID_negPS10G_1_A => return "L1PHID_negPS10G_1_A";
       when L6PHIA_neg2S_3_A => return "L6PHIA_neg2S_3_A";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_AS_36) return string is
  begin
    case val is
       when L4PHIDn2 => return "L4PHIDn2";
       when L3PHICn6 => return "L3PHICn6";
       when L5PHIBn1 => return "L5PHIBn1";
       when L3PHIDn1 => return "L3PHIDn1";
       when L1PHIHn3 => return "L1PHIHn3";
       when L1PHIBn1 => return "L1PHIBn1";
       when L1PHIAn1 => return "L1PHIAn1";
       when L2PHICn6 => return "L2PHICn6";
       when L1PHIGn3 => return "L1PHIGn3";
       when L4PHIAn3 => return "L4PHIAn3";
       when L2PHICn4 => return "L2PHICn4";
       when L2PHICn2 => return "L2PHICn2";
       when L1PHIDn2 => return "L1PHIDn2";
       when L3PHICn2 => return "L3PHICn2";
       when L4PHIBn4 => return "L4PHIBn4";
       when L2PHIDn4 => return "L2PHIDn4";
       when L4PHIBn1 => return "L4PHIBn1";
       when L5PHIAn2 => return "L5PHIAn2";
       when L1PHIDn1 => return "L1PHIDn1";
       when L4PHIDn1 => return "L4PHIDn1";
       when L1PHICn3 => return "L1PHICn3";
       when L1PHICn4 => return "L1PHICn4";
       when L1PHIGn2 => return "L1PHIGn2";
       when L2PHIBn3 => return "L2PHIBn3";
       when L3PHIBn2 => return "L3PHIBn2";
       when L3PHICn4 => return "L3PHICn4";
       when L1PHIEn1 => return "L1PHIEn1";
       when L6PHIDn3 => return "L6PHIDn3";
       when L1PHIFn3 => return "L1PHIFn3";
       when L1PHIAn3 => return "L1PHIAn3";
       when L2PHICn7 => return "L2PHICn7";
       when L6PHICn2 => return "L6PHICn2";
       when L2PHIBn6 => return "L2PHIBn6";
       when L5PHIBn3 => return "L5PHIBn3";
       when L2PHICn1 => return "L2PHICn1";
       when L3PHIDn3 => return "L3PHIDn3";
       when L4PHICn4 => return "L4PHICn4";
       when L1PHIBn2 => return "L1PHIBn2";
       when L4PHIAn2 => return "L4PHIAn2";
       when L2PHIBn1 => return "L2PHIBn1";
       when L5PHIDn2 => return "L5PHIDn2";
       when L2PHIAn6 => return "L2PHIAn6";
       when L3PHIDn2 => return "L3PHIDn2";
       when L2PHIBn7 => return "L2PHIBn7";
       when L3PHIBn6 => return "L3PHIBn6";
       when L2PHICn5 => return "L2PHICn5";
       when L2PHIAn1 => return "L2PHIAn1";
       when L2PHIBn8 => return "L2PHIBn8";
       when L2PHIBn5 => return "L2PHIBn5";
       when L6PHIBn3 => return "L6PHIBn3";
       when L1PHIFn1 => return "L1PHIFn1";
       when L6PHIAn2 => return "L6PHIAn2";
       when L6PHIDn2 => return "L6PHIDn2";
       when L5PHICn1 => return "L5PHICn1";
       when L5PHIDn1 => return "L5PHIDn1";
       when L1PHIHn2 => return "L1PHIHn2";
       when L1PHIEn3 => return "L1PHIEn3";
       when L4PHIBn3 => return "L4PHIBn3";
       when L4PHIAn1 => return "L4PHIAn1";
       when L5PHICn3 => return "L5PHICn3";
       when L4PHIBn2 => return "L4PHIBn2";
       when L3PHIBn5 => return "L3PHIBn5";
       when L3PHIBn4 => return "L3PHIBn4";
       when L3PHICn3 => return "L3PHICn3";
       when L1PHIFn4 => return "L1PHIFn4";
       when L6PHICn1 => return "L6PHICn1";
       when L2PHIAn5 => return "L2PHIAn5";
       when L3PHIBn3 => return "L3PHIBn3";
       when L3PHICn1 => return "L3PHICn1";
       when L2PHIBn2 => return "L2PHIBn2";
       when L5PHIBn2 => return "L5PHIBn2";
       when L6PHIBn2 => return "L6PHIBn2";
       when L4PHIDn3 => return "L4PHIDn3";
       when L1PHICn2 => return "L1PHICn2";
       when L6PHICn3 => return "L6PHICn3";
       when L6PHICn4 => return "L6PHICn4";
       when L2PHICn3 => return "L2PHICn3";
       when L1PHIFn2 => return "L1PHIFn2";
       when L4PHICn3 => return "L4PHICn3";
       when L2PHIDn2 => return "L2PHIDn2";
       when L3PHIDn4 => return "L3PHIDn4";
       when L1PHIGn1 => return "L1PHIGn1";
       when L6PHIDn1 => return "L6PHIDn1";
       when L2PHIAn3 => return "L2PHIAn3";
       when L6PHIBn1 => return "L6PHIBn1";
       when L1PHIHn1 => return "L1PHIHn1";
       when L2PHIAn4 => return "L2PHIAn4";
       when L2PHIDn3 => return "L2PHIDn3";
       when L3PHIAn2 => return "L3PHIAn2";
       when L1PHIAn2 => return "L1PHIAn2";
       when L3PHIBn1 => return "L3PHIBn1";
       when L2PHIDn1 => return "L2PHIDn1";
       when L5PHIAn1 => return "L5PHIAn1";
       when L2PHIAn2 => return "L2PHIAn2";
       when L6PHIAn3 => return "L6PHIAn3";
       when L1PHICn1 => return "L1PHICn1";
       when L2PHIBn4 => return "L2PHIBn4";
       when L4PHICn2 => return "L4PHICn2";
       when L6PHIBn4 => return "L6PHIBn4";
       when L3PHIAn3 => return "L3PHIAn3";
       when L1PHIDn3 => return "L1PHIDn3";
       when L1PHIBn3 => return "L1PHIBn3";
       when L4PHICn1 => return "L4PHICn1";
       when L6PHIAn1 => return "L6PHIAn1";
       when L2PHIDn6 => return "L2PHIDn6";
       when L3PHICn5 => return "L3PHICn5";
       when L2PHIDn5 => return "L2PHIDn5";
       when L5PHICn2 => return "L5PHICn2";
       when L3PHIAn1 => return "L3PHIAn1";
       when L1PHIEn2 => return "L1PHIEn2";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSME_17) return string is
  begin
    case val is
       when L5PHID28n1 => return "L5PHID28n1";
       when L5PHIC23n1 => return "L5PHIC23n1";
       when L4PHIB15n1 => return "L4PHIB15n1";
       when L4PHIC21n1 => return "L4PHIC21n1";
       when L4PHIA4n1 => return "L4PHIA4n1";
       when L5PHID25n1 => return "L5PHID25n1";
       when L6PHIB12n1 => return "L6PHIB12n1";
       when L6PHIC18n1 => return "L6PHIC18n1";
       when L4PHIB14n1 => return "L4PHIB14n1";
       when L4PHIA3n1 => return "L4PHIA3n1";
       when L4PHIB10n1 => return "L4PHIB10n1";
       when L5PHIB13n1 => return "L5PHIB13n1";
       when L6PHIB9n1 => return "L6PHIB9n1";
       when L6PHID32n1 => return "L6PHID32n1";
       when L5PHIA5n1 => return "L5PHIA5n1";
       when L5PHIA1n1 => return "L5PHIA1n1";
       when L4PHID28n1 => return "L4PHID28n1";
       when L5PHIC17n1 => return "L5PHIC17n1";
       when L4PHID25n1 => return "L4PHID25n1";
       when L4PHIC22n1 => return "L4PHIC22n1";
       when L6PHIA2n1 => return "L6PHIA2n1";
       when L6PHIA6n1 => return "L6PHIA6n1";
       when L4PHIA7n1 => return "L4PHIA7n1";
       when L6PHIC21n1 => return "L6PHIC21n1";
       when L5PHIC22n1 => return "L5PHIC22n1";
       when L4PHIB9n1 => return "L4PHIB9n1";
       when L4PHID30n1 => return "L4PHID30n1";
       when L5PHIB14n1 => return "L5PHIB14n1";
       when L6PHIB16n1 => return "L6PHIB16n1";
       when L6PHID26n1 => return "L6PHID26n1";
       when L6PHIA3n1 => return "L6PHIA3n1";
       when L6PHIC17n1 => return "L6PHIC17n1";
       when L5PHID31n1 => return "L5PHID31n1";
       when L6PHIC22n1 => return "L6PHIC22n1";
       when L6PHID30n1 => return "L6PHID30n1";
       when L6PHID31n1 => return "L6PHID31n1";
       when L5PHIB15n1 => return "L5PHIB15n1";
       when L4PHIC24n1 => return "L4PHIC24n1";
       when L5PHID32n1 => return "L5PHID32n1";
       when L4PHIC17n1 => return "L4PHIC17n1";
       when L4PHID29n1 => return "L4PHID29n1";
       when L4PHIA6n1 => return "L4PHIA6n1";
       when L4PHID27n1 => return "L4PHID27n1";
       when L6PHIB13n1 => return "L6PHIB13n1";
       when L6PHIC24n1 => return "L6PHIC24n1";
       when L5PHIB11n1 => return "L5PHIB11n1";
       when L5PHID26n1 => return "L5PHID26n1";
       when L4PHIC20n1 => return "L4PHIC20n1";
       when L5PHIC24n1 => return "L5PHIC24n1";
       when L5PHIA2n1 => return "L5PHIA2n1";
       when L5PHID30n1 => return "L5PHID30n1";
       when L5PHIB10n1 => return "L5PHIB10n1";
       when L6PHIC19n1 => return "L6PHIC19n1";
       when L5PHIA6n1 => return "L5PHIA6n1";
       when L4PHID31n1 => return "L4PHID31n1";
       when L5PHID29n1 => return "L5PHID29n1";
       when L5PHIA8n1 => return "L5PHIA8n1";
       when L4PHIA8n1 => return "L4PHIA8n1";
       when L4PHIB16n1 => return "L4PHIB16n1";
       when L4PHID32n1 => return "L4PHID32n1";
       when L6PHIB11n1 => return "L6PHIB11n1";
       when L5PHIC20n1 => return "L5PHIC20n1";
       when L4PHID26n1 => return "L4PHID26n1";
       when L4PHIB13n1 => return "L4PHIB13n1";
       when L6PHIC23n1 => return "L6PHIC23n1";
       when L6PHIA8n1 => return "L6PHIA8n1";
       when L4PHIA2n1 => return "L4PHIA2n1";
       when L5PHID27n1 => return "L5PHID27n1";
       when L6PHIA4n1 => return "L6PHIA4n1";
       when L5PHIB16n1 => return "L5PHIB16n1";
       when L5PHIC21n1 => return "L5PHIC21n1";
       when L5PHIC19n1 => return "L5PHIC19n1";
       when L6PHIB10n1 => return "L6PHIB10n1";
       when L6PHIB15n1 => return "L6PHIB15n1";
       when L6PHIB14n1 => return "L6PHIB14n1";
       when L5PHIA3n1 => return "L5PHIA3n1";
       when L5PHIA4n1 => return "L5PHIA4n1";
       when L5PHIB12n1 => return "L5PHIB12n1";
       when L4PHIB11n1 => return "L4PHIB11n1";
       when L6PHID28n1 => return "L6PHID28n1";
       when L4PHIB12n1 => return "L4PHIB12n1";
       when L5PHIC18n1 => return "L5PHIC18n1";
       when L4PHIC19n1 => return "L4PHIC19n1";
       when L6PHIA7n1 => return "L6PHIA7n1";
       when L4PHIA1n1 => return "L4PHIA1n1";
       when L6PHIA5n1 => return "L6PHIA5n1";
       when L6PHID29n1 => return "L6PHID29n1";
       when L4PHIC18n1 => return "L4PHIC18n1";
       when L5PHIB9n1 => return "L5PHIB9n1";
       when L4PHIC23n1 => return "L4PHIC23n1";
       when L6PHID27n1 => return "L6PHID27n1";
       when L6PHID25n1 => return "L6PHID25n1";
       when L6PHIC20n1 => return "L6PHIC20n1";
       when L5PHIA7n1 => return "L5PHIA7n1";
       when L4PHIA5n1 => return "L4PHIA5n1";
       when L6PHIA1n1 => return "L6PHIA1n1";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSME_16) return string is
  begin
    case val is
       when L2PHIC21n1 => return "L2PHIC21n1";
       when L2PHID31n1 => return "L2PHID31n1";
       when L2PHIB10n1 => return "L2PHIB10n1";
       when L1PHIF22n1 => return "L1PHIF22n1";
       when L3PHID25n1 => return "L3PHID25n1";
       when L1PHIA2n1 => return "L1PHIA2n1";
       when L1PHID15n1 => return "L1PHID15n1";
       when L1PHIA3n1 => return "L1PHIA3n1";
       when L3PHIA3n1 => return "L3PHIA3n1";
       when L3PHIC23n1 => return "L3PHIC23n1";
       when L1PHID16n1 => return "L1PHID16n1";
       when L1PHIE17n1 => return "L1PHIE17n1";
       when L3PHID26n1 => return "L3PHID26n1";
       when L2PHID29n1 => return "L2PHID29n1";
       when L2PHID30n1 => return "L2PHID30n1";
       when L2PHIA4n1 => return "L2PHIA4n1";
       when L1PHIG28n1 => return "L1PHIG28n1";
       when L2PHIC19n1 => return "L2PHIC19n1";
       when L1PHIA4n1 => return "L1PHIA4n1";
       when L1PHIC9n1 => return "L1PHIC9n1";
       when L3PHIB11n1 => return "L3PHIB11n1";
       when L1PHIF21n1 => return "L1PHIF21n1";
       when L1PHIF23n1 => return "L1PHIF23n1";
       when L1PHIE19n1 => return "L1PHIE19n1";
       when L2PHIC24n1 => return "L2PHIC24n1";
       when L2PHIB9n1 => return "L2PHIB9n1";
       when L3PHIC21n1 => return "L3PHIC21n1";
       when L3PHIA5n1 => return "L3PHIA5n1";
       when L3PHIB10n1 => return "L3PHIB10n1";
       when L3PHID28n1 => return "L3PHID28n1";
       when L3PHID32n1 => return "L3PHID32n1";
       when L3PHID30n1 => return "L3PHID30n1";
       when L2PHIB14n1 => return "L2PHIB14n1";
       when L2PHIC17n1 => return "L2PHIC17n1";
       when L1PHIH30n1 => return "L1PHIH30n1";
       when L1PHIG25n1 => return "L1PHIG25n1";
       when L1PHIH31n1 => return "L1PHIH31n1";
       when L3PHIA4n1 => return "L3PHIA4n1";
       when L3PHIA7n1 => return "L3PHIA7n1";
       when L2PHIB16n1 => return "L2PHIB16n1";
       when L3PHIC17n1 => return "L3PHIC17n1";
       when L1PHIH32n1 => return "L1PHIH32n1";
       when L2PHIC18n1 => return "L2PHIC18n1";
       when L2PHIA7n1 => return "L2PHIA7n1";
       when L3PHIA6n1 => return "L3PHIA6n1";
       when L3PHIA8n1 => return "L3PHIA8n1";
       when L3PHIB9n1 => return "L3PHIB9n1";
       when L2PHID32n1 => return "L2PHID32n1";
       when L3PHIC22n1 => return "L3PHIC22n1";
       when L1PHIC10n1 => return "L1PHIC10n1";
       when L2PHIA5n1 => return "L2PHIA5n1";
       when L2PHIC23n1 => return "L2PHIC23n1";
       when L1PHIA1n1 => return "L1PHIA1n1";
       when L1PHIC12n1 => return "L1PHIC12n1";
       when L1PHIC11n1 => return "L1PHIC11n1";
       when L1PHID13n1 => return "L1PHID13n1";
       when L2PHIC20n1 => return "L2PHIC20n1";
       when L2PHIA6n1 => return "L2PHIA6n1";
       when L3PHIC18n1 => return "L3PHIC18n1";
       when L1PHIE20n1 => return "L1PHIE20n1";
       when L2PHIA3n1 => return "L2PHIA3n1";
       when L3PHIB14n1 => return "L3PHIB14n1";
       when L2PHIA8n1 => return "L2PHIA8n1";
       when L1PHIB7n1 => return "L1PHIB7n1";
       when L1PHIB5n1 => return "L1PHIB5n1";
       when L1PHIB8n1 => return "L1PHIB8n1";
       when L2PHID26n1 => return "L2PHID26n1";
       when L1PHIG26n1 => return "L1PHIG26n1";
       when L2PHIB13n1 => return "L2PHIB13n1";
       when L2PHIB15n1 => return "L2PHIB15n1";
       when L2PHID28n1 => return "L2PHID28n1";
       when L3PHID29n1 => return "L3PHID29n1";
       when L1PHID14n1 => return "L1PHID14n1";
       when L1PHIB6n1 => return "L1PHIB6n1";
       when L2PHIA2n1 => return "L2PHIA2n1";
       when L3PHIB15n1 => return "L3PHIB15n1";
       when L3PHID31n1 => return "L3PHID31n1";
       when L3PHIC24n1 => return "L3PHIC24n1";
       when L2PHIA1n1 => return "L2PHIA1n1";
       when L3PHIA1n1 => return "L3PHIA1n1";
       when L3PHIC19n1 => return "L3PHIC19n1";
       when L1PHIE18n1 => return "L1PHIE18n1";
       when L1PHIG27n1 => return "L1PHIG27n1";
       when L3PHIB16n1 => return "L3PHIB16n1";
       when L3PHIB13n1 => return "L3PHIB13n1";
       when L2PHIB11n1 => return "L2PHIB11n1";
       when L2PHIB12n1 => return "L2PHIB12n1";
       when L1PHIH29n1 => return "L1PHIH29n1";
       when L2PHID25n1 => return "L2PHID25n1";
       when L2PHID27n1 => return "L2PHID27n1";
       when L1PHIF24n1 => return "L1PHIF24n1";
       when L3PHID27n1 => return "L3PHID27n1";
       when L3PHIB12n1 => return "L3PHIB12n1";
       when L3PHIC20n1 => return "L3PHIC20n1";
       when L2PHIC22n1 => return "L2PHIC22n1";
       when L3PHIA2n1 => return "L3PHIA2n1";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSTE_22) return string is
  begin
    case val is
       when L2PHIJ6n3 => return "L2PHIJ6n3";
       when L3PHID15n2 => return "L3PHID15n2";
       when L2PHIJ6n2 => return "L2PHIJ6n2";
       when L3PHID13n5 => return "L3PHID13n5";
       when L1PHIA2n3 => return "L1PHIA2n3";
       when L1PHIB6n2 => return "L1PHIB6n2";
       when L1PHIB8n3 => return "L1PHIB8n3";
       when L1PHIA4n2 => return "L1PHIA4n2";
       when L3PHID14n3 => return "L3PHID14n3";
       when L1PHIE19n3 => return "L1PHIE19n3";
       when L2PHIK10n2 => return "L2PHIK10n2";
       when L1PHIB6n3 => return "L1PHIB6n3";
       when L1PHIE17n4 => return "L1PHIE17n4";
       when L1PHID16n3 => return "L1PHID16n3";
       when L3PHIC9n5 => return "L3PHIC9n5";
       when L1PHIG25n3 => return "L1PHIG25n3";
       when L3PHID16n3 => return "L3PHID16n3";
       when L1PHID16n4 => return "L1PHID16n4";
       when L2PHIK12n1 => return "L2PHIK12n1";
       when L1PHIA1n3 => return "L1PHIA1n3";
       when L1PHIF23n2 => return "L1PHIF23n2";
       when L1PHIH31n4 => return "L1PHIH31n4";
       when L1PHIC12n1 => return "L1PHIC12n1";
       when L1PHIG25n2 => return "L1PHIG25n2";
       when L1PHIG26n3 => return "L1PHIG26n3";
       when L1PHIB7n1 => return "L1PHIB7n1";
       when L3PHIA2n4 => return "L3PHIA2n4";
       when L3PHIA2n5 => return "L3PHIA2n5";
       when L2PHII3n3 => return "L2PHII3n3";
       when L1PHIF21n4 => return "L1PHIF21n4";
       when L1PHIB8n2 => return "L1PHIB8n2";
       when L3PHIA3n1 => return "L3PHIA3n1";
       when L1PHIH32n2 => return "L1PHIH32n2";
       when L3PHIC10n6 => return "L3PHIC10n6";
       when L3PHIC11n6 => return "L3PHIC11n6";
       when L2PHIL13n1 => return "L2PHIL13n1";
       when L2PHIL15n3 => return "L2PHIL15n3";
       when L3PHIB5n3 => return "L3PHIB5n3";
       when L2PHIJ8n1 => return "L2PHIJ8n1";
       when L1PHIH32n3 => return "L1PHIH32n3";
       when L1PHIF24n2 => return "L1PHIF24n2";
       when L1PHIA1n2 => return "L1PHIA1n2";
       when L1PHIF23n5 => return "L1PHIF23n5";
       when L2PHIJ8n3 => return "L2PHIJ8n3";
       when L1PHIG27n2 => return "L1PHIG27n2";
       when L1PHIG26n2 => return "L1PHIG26n2";
       when L1PHIA4n1 => return "L1PHIA4n1";
       when L3PHID16n2 => return "L3PHID16n2";
       when L1PHIB6n5 => return "L1PHIB6n5";
       when L3PHIA1n4 => return "L3PHIA1n4";
       when L2PHIL16n1 => return "L2PHIL16n1";
       when L1PHIG28n2 => return "L1PHIG28n2";
       when L2PHIL13n3 => return "L2PHIL13n3";
       when L3PHIA4n1 => return "L3PHIA4n1";
       when L3PHID14n5 => return "L3PHID14n5";
       when L1PHIG27n4 => return "L1PHIG27n4";
       when L2PHIK12n2 => return "L2PHIK12n2";
       when L1PHIC11n4 => return "L1PHIC11n4";
       when L3PHIC11n5 => return "L3PHIC11n5";
       when L3PHIB6n2 => return "L3PHIB6n2";
       when L1PHIB5n2 => return "L1PHIB5n2";
       when L3PHIC9n6 => return "L3PHIC9n6";
       when L1PHIC11n1 => return "L1PHIC11n1";
       when L1PHIF22n1 => return "L1PHIF22n1";
       when L1PHIC11n2 => return "L1PHIC11n2";
       when L3PHID15n1 => return "L3PHID15n1";
       when L1PHIG27n5 => return "L1PHIG27n5";
       when L3PHID15n3 => return "L3PHID15n3";
       when L1PHIE17n3 => return "L1PHIE17n3";
       when L1PHIC12n3 => return "L1PHIC12n3";
       when L1PHIB5n1 => return "L1PHIB5n1";
       when L1PHIC10n4 => return "L1PHIC10n4";
       when L1PHID14n2 => return "L1PHID14n2";
       when L1PHIC9n3 => return "L1PHIC9n3";
       when L3PHIB6n5 => return "L3PHIB6n5";
       when L1PHIH29n1 => return "L1PHIH29n1";
       when L1PHID14n4 => return "L1PHID14n4";
       when L1PHIE17n5 => return "L1PHIE17n5";
       when L1PHIB8n1 => return "L1PHIB8n1";
       when L1PHIE20n4 => return "L1PHIE20n4";
       when L1PHIG28n1 => return "L1PHIG28n1";
       when L3PHIC12n4 => return "L3PHIC12n4";
       when L1PHIA3n4 => return "L1PHIA3n4";
       when L1PHID15n1 => return "L1PHID15n1";
       when L1PHIE17n1 => return "L1PHIE17n1";
       when L3PHIB5n5 => return "L3PHIB5n5";
       when L1PHIG25n4 => return "L1PHIG25n4";
       when L3PHID16n4 => return "L3PHID16n4";
       when L1PHIE20n3 => return "L1PHIE20n3";
       when L1PHID16n2 => return "L1PHID16n2";
       when L3PHIC12n5 => return "L3PHIC12n5";
       when L2PHIK11n2 => return "L2PHIK11n2";
       when L3PHID13n3 => return "L3PHID13n3";
       when L3PHIB7n2 => return "L3PHIB7n2";
       when L1PHIF23n4 => return "L1PHIF23n4";
       when L1PHIC10n5 => return "L1PHIC10n5";
       when L3PHID13n2 => return "L3PHID13n2";
       when L2PHII4n1 => return "L2PHII4n1";
       when L3PHIB6n4 => return "L3PHIB6n4";
       when L2PHII3n1 => return "L2PHII3n1";
       when L2PHII1n2 => return "L2PHII1n2";
       when L2PHIL14n1 => return "L2PHIL14n1";
       when L1PHIA4n4 => return "L1PHIA4n4";
       when L1PHIE18n1 => return "L1PHIE18n1";
       when L3PHIA3n2 => return "L3PHIA3n2";
       when L2PHIK9n3 => return "L2PHIK9n3";
       when L3PHIC11n1 => return "L3PHIC11n1";
       when L2PHII3n2 => return "L2PHII3n2";
       when L1PHIE18n2 => return "L1PHIE18n2";
       when L1PHIH32n1 => return "L1PHIH32n1";
       when L1PHID13n2 => return "L1PHID13n2";
       when L3PHIC10n3 => return "L3PHIC10n3";
       when L1PHIH30n4 => return "L1PHIH30n4";
       when L1PHIA3n2 => return "L1PHIA3n2";
       when L1PHIE17n2 => return "L1PHIE17n2";
       when L1PHIB6n1 => return "L1PHIB6n1";
       when L3PHID14n4 => return "L3PHID14n4";
       when L2PHIK10n1 => return "L2PHIK10n1";
       when L1PHIF24n5 => return "L1PHIF24n5";
       when L2PHII4n3 => return "L2PHII4n3";
       when L2PHIK9n1 => return "L2PHIK9n1";
       when L2PHIJ7n2 => return "L2PHIJ7n2";
       when L3PHIB7n4 => return "L3PHIB7n4";
       when L3PHID13n1 => return "L3PHID13n1";
       when L3PHIC12n3 => return "L3PHIC12n3";
       when L1PHIC10n1 => return "L1PHIC10n1";
       when L3PHIB8n2 => return "L3PHIB8n2";
       when L2PHIJ5n1 => return "L2PHIJ5n1";
       when L2PHIJ6n1 => return "L2PHIJ6n1";
       when L1PHIF21n1 => return "L1PHIF21n1";
       when L1PHIF21n3 => return "L1PHIF21n3";
       when L1PHIC9n5 => return "L1PHIC9n5";
       when L1PHIF22n2 => return "L1PHIF22n2";
       when L1PHIC12n2 => return "L1PHIC12n2";
       when L1PHIH31n1 => return "L1PHIH31n1";
       when L1PHIG25n5 => return "L1PHIG25n5";
       when L1PHIB7n4 => return "L1PHIB7n4";
       when L1PHIA4n3 => return "L1PHIA4n3";
       when L3PHIB5n4 => return "L3PHIB5n4";
       when L1PHID13n1 => return "L1PHID13n1";
       when L1PHIF24n3 => return "L1PHIF24n3";
       when L1PHIG28n5 => return "L1PHIG28n5";
       when L1PHIE18n4 => return "L1PHIE18n4";
       when L3PHIB7n3 => return "L3PHIB7n3";
       when L2PHIL14n2 => return "L2PHIL14n2";
       when L2PHIK11n3 => return "L2PHIK11n3";
       when L3PHIC9n2 => return "L3PHIC9n2";
       when L3PHIC11n3 => return "L3PHIC11n3";
       when L3PHIB7n1 => return "L3PHIB7n1";
       when L1PHIE19n2 => return "L1PHIE19n2";
       when L3PHIA4n3 => return "L3PHIA4n3";
       when L1PHID13n4 => return "L1PHID13n4";
       when L1PHIF24n4 => return "L1PHIF24n4";
       when L2PHIK12n3 => return "L2PHIK12n3";
       when L3PHIB8n4 => return "L3PHIB8n4";
       when L3PHIB7n6 => return "L3PHIB7n6";
       when L1PHIH30n5 => return "L1PHIH30n5";
       when L2PHIJ8n2 => return "L2PHIJ8n2";
       when L1PHIC11n3 => return "L1PHIC11n3";
       when L1PHIH30n1 => return "L1PHIH30n1";
       when L3PHIC10n5 => return "L3PHIC10n5";
       when L3PHID15n6 => return "L3PHID15n6";
       when L1PHIC10n2 => return "L1PHIC10n2";
       when L1PHIC10n3 => return "L1PHIC10n3";
       when L3PHID16n1 => return "L3PHID16n1";
       when L1PHIG28n4 => return "L1PHIG28n4";
       when L1PHID13n5 => return "L1PHID13n5";
       when L1PHIG28n3 => return "L1PHIG28n3";
       when L3PHIC9n1 => return "L3PHIC9n1";
       when L1PHID15n5 => return "L1PHID15n5";
       when L1PHIH29n2 => return "L1PHIH29n2";
       when L3PHIA3n3 => return "L3PHIA3n3";
       when L1PHIH30n3 => return "L1PHIH30n3";
       when L3PHIA3n4 => return "L3PHIA3n4";
       when L1PHIA4n5 => return "L1PHIA4n5";
       when L1PHIF22n3 => return "L1PHIF22n3";
       when L1PHID14n5 => return "L1PHID14n5";
       when L3PHIA3n5 => return "L3PHIA3n5";
       when L1PHIA3n5 => return "L1PHIA3n5";
       when L1PHIH31n3 => return "L1PHIH31n3";
       when L2PHIJ5n2 => return "L2PHIJ5n2";
       when L1PHIB7n5 => return "L1PHIB7n5";
       when L2PHIL15n1 => return "L2PHIL15n1";
       when L1PHIA3n1 => return "L1PHIA3n1";
       when L1PHIF22n5 => return "L1PHIF22n5";
       when L2PHIL14n3 => return "L2PHIL14n3";
       when L2PHII2n1 => return "L2PHII2n1";
       when L1PHID15n3 => return "L1PHID15n3";
       when L1PHIG27n1 => return "L1PHIG27n1";
       when L3PHIC12n2 => return "L3PHIC12n2";
       when L1PHIC12n4 => return "L1PHIC12n4";
       when L3PHIA2n1 => return "L3PHIA2n1";
       when L1PHIB5n3 => return "L1PHIB5n3";
       when L3PHIA1n2 => return "L3PHIA1n2";
       when L3PHIC11n4 => return "L3PHIC11n4";
       when L1PHIF23n3 => return "L1PHIF23n3";
       when L1PHIH30n2 => return "L1PHIH30n2";
       when L1PHIF21n5 => return "L1PHIF21n5";
       when L1PHIA2n4 => return "L1PHIA2n4";
       when L3PHIC12n6 => return "L3PHIC12n6";
       when L3PHIB5n2 => return "L3PHIB5n2";
       when L3PHIA1n3 => return "L3PHIA1n3";
       when L1PHIH29n5 => return "L1PHIH29n5";
       when L1PHIB5n5 => return "L1PHIB5n5";
       when L3PHIB7n5 => return "L3PHIB7n5";
       when L3PHIA4n6 => return "L3PHIA4n6";
       when L1PHIF21n2 => return "L1PHIF21n2";
       when L3PHIA2n2 => return "L3PHIA2n2";
       when L1PHIH31n2 => return "L1PHIH31n2";
       when L1PHIF24n1 => return "L1PHIF24n1";
       when L1PHIC9n2 => return "L1PHIC9n2";
       when L3PHIC9n4 => return "L3PHIC9n4";
       when L3PHIA1n1 => return "L3PHIA1n1";
       when L3PHID13n6 => return "L3PHID13n6";
       when L3PHIC12n1 => return "L3PHIC12n1";
       when L1PHIA2n1 => return "L1PHIA2n1";
       when L1PHIB8n5 => return "L1PHIB8n5";
       when L3PHIA3n6 => return "L3PHIA3n6";
       when L3PHID14n2 => return "L3PHID14n2";
       when L1PHIC12n5 => return "L1PHIC12n5";
       when L2PHII1n1 => return "L2PHII1n1";
       when L2PHIJ5n3 => return "L2PHIJ5n3";
       when L1PHIB6n4 => return "L1PHIB6n4";
       when L3PHIB5n6 => return "L3PHIB5n6";
       when L3PHIC11n2 => return "L3PHIC11n2";
       when L1PHIF22n4 => return "L1PHIF22n4";
       when L2PHII2n2 => return "L2PHII2n2";
       when L2PHIL16n2 => return "L2PHIL16n2";
       when L1PHIB7n2 => return "L1PHIB7n2";
       when L2PHIK9n2 => return "L2PHIK9n2";
       when L3PHIA4n4 => return "L3PHIA4n4";
       when L2PHIL13n2 => return "L2PHIL13n2";
       when L3PHIC10n2 => return "L3PHIC10n2";
       when L3PHIB8n1 => return "L3PHIB8n1";
       when L1PHIA3n3 => return "L1PHIA3n3";
       when L3PHIC10n1 => return "L3PHIC10n1";
       when L3PHID15n4 => return "L3PHID15n4";
       when L1PHIE20n5 => return "L1PHIE20n5";
       when L1PHID13n3 => return "L1PHID13n3";
       when L1PHIE18n5 => return "L1PHIE18n5";
       when L2PHIL15n2 => return "L2PHIL15n2";
       when L1PHIE20n1 => return "L1PHIE20n1";
       when L1PHID16n5 => return "L1PHID16n5";
       when L3PHID15n5 => return "L3PHID15n5";
       when L3PHIB6n3 => return "L3PHIB6n3";
       when L3PHID14n6 => return "L3PHID14n6";
       when L1PHIB7n3 => return "L1PHIB7n3";
       when L3PHIB6n6 => return "L3PHIB6n6";
       when L1PHIA1n1 => return "L1PHIA1n1";
       when L1PHIE19n4 => return "L1PHIE19n4";
       when L1PHIH29n3 => return "L1PHIH29n3";
       when L1PHID14n3 => return "L1PHID14n3";
       when L1PHIE19n1 => return "L1PHIE19n1";
       when L1PHIB8n4 => return "L1PHIB8n4";
       when L3PHID14n1 => return "L3PHID14n1";
       when L1PHIG26n4 => return "L1PHIG26n4";
       when L1PHIE19n5 => return "L1PHIE19n5";
       when L1PHIA2n2 => return "L1PHIA2n2";
       when L2PHIK11n1 => return "L2PHIK11n1";
       when L3PHIC10n4 => return "L3PHIC10n4";
       when L1PHID16n1 => return "L1PHID16n1";
       when L3PHIA2n3 => return "L3PHIA2n3";
       when L3PHIB8n6 => return "L3PHIB8n6";
       when L1PHIC11n5 => return "L1PHIC11n5";
       when L1PHIE20n2 => return "L1PHIE20n2";
       when L3PHIA4n2 => return "L3PHIA4n2";
       when L1PHID14n1 => return "L1PHID14n1";
       when L2PHII2n3 => return "L2PHII2n3";
       when L3PHIB5n1 => return "L3PHIB5n1";
       when L2PHIK10n3 => return "L2PHIK10n3";
       when L1PHIE18n3 => return "L1PHIE18n3";
       when L1PHIC9n1 => return "L1PHIC9n1";
       when L3PHID13n4 => return "L3PHID13n4";
       when L3PHIA2n6 => return "L3PHIA2n6";
       when L2PHIJ7n3 => return "L2PHIJ7n3";
       when L2PHIJ7n1 => return "L2PHIJ7n1";
       when L1PHIC9n4 => return "L1PHIC9n4";
       when L1PHIG26n1 => return "L1PHIG26n1";
       when L3PHIB6n1 => return "L3PHIB6n1";
       when L1PHIG27n3 => return "L1PHIG27n3";
       when L1PHID15n2 => return "L1PHID15n2";
       when L1PHIG26n5 => return "L1PHIG26n5";
       when L1PHID15n4 => return "L1PHID15n4";
       when L3PHIB8n5 => return "L3PHIB8n5";
       when L1PHIF23n1 => return "L1PHIF23n1";
       when L3PHIB8n3 => return "L3PHIB8n3";
       when L2PHII4n2 => return "L2PHII4n2";
       when L3PHIA4n5 => return "L3PHIA4n5";
       when L1PHIG25n1 => return "L1PHIG25n1";
       when L1PHIB5n4 => return "L1PHIB5n4";
       when L1PHIH29n4 => return "L1PHIH29n4";
       when L3PHIC9n3 => return "L3PHIC9n3";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSTE_17) return string is
  begin
    case val is
       when L6PHIC22n1 => return "L6PHIC22n1";
       when L6PHID27n1 => return "L6PHID27n1";
       when L6PHID26n1 => return "L6PHID26n1";
       when L6PHIC24n2 => return "L6PHIC24n2";
       when L6PHIB11n4 => return "L6PHIB11n4";
       when L6PHIA6n3 => return "L6PHIA6n3";
       when L6PHIB13n2 => return "L6PHIB13n2";
       when L6PHIA8n3 => return "L6PHIA8n3";
       when L6PHID25n1 => return "L6PHID25n1";
       when L6PHIB15n3 => return "L6PHIB15n3";
       when L6PHID29n1 => return "L6PHID29n1";
       when L6PHIB14n3 => return "L6PHIB14n3";
       when L4PHID25n2 => return "L4PHID25n2";
       when L6PHIB12n1 => return "L6PHIB12n1";
       when L4PHIA4n1 => return "L4PHIA4n1";
       when L6PHIB15n1 => return "L6PHIB15n1";
       when L4PHIA6n1 => return "L4PHIA6n1";
       when L6PHID25n3 => return "L6PHID25n3";
       when L6PHID27n4 => return "L6PHID27n4";
       when L6PHIC17n3 => return "L6PHIC17n3";
       when L4PHIC18n1 => return "L4PHIC18n1";
       when L6PHID25n2 => return "L6PHID25n2";
       when L6PHIB12n4 => return "L6PHIB12n4";
       when L6PHID28n1 => return "L6PHID28n1";
       when L6PHIC19n1 => return "L6PHIC19n1";
       when L4PHIC22n2 => return "L4PHIC22n2";
       when L6PHID29n4 => return "L6PHID29n4";
       when L6PHIC19n2 => return "L6PHIC19n2";
       when L6PHIB14n2 => return "L6PHIB14n2";
       when L6PHIB11n1 => return "L6PHIB11n1";
       when L6PHIC18n1 => return "L6PHIC18n1";
       when L6PHIB9n2 => return "L6PHIB9n2";
       when L4PHIC20n2 => return "L4PHIC20n2";
       when L6PHIB10n3 => return "L6PHIB10n3";
       when L4PHIC18n3 => return "L4PHIC18n3";
       when L4PHIB13n3 => return "L4PHIB13n3";
       when L4PHIB14n3 => return "L4PHIB14n3";
       when L4PHIB14n2 => return "L4PHIB14n2";
       when L4PHIB13n2 => return "L4PHIB13n2";
       when L4PHIB16n2 => return "L4PHIB16n2";
       when L6PHIA3n3 => return "L6PHIA3n3";
       when L4PHIC17n3 => return "L4PHIC17n3";
       when L6PHID27n2 => return "L6PHID27n2";
       when L6PHIB11n3 => return "L6PHIB11n3";
       when L6PHIB12n2 => return "L6PHIB12n2";
       when L6PHID28n2 => return "L6PHID28n2";
       when L6PHIA7n3 => return "L6PHIA7n3";
       when L4PHID25n1 => return "L4PHID25n1";
       when L4PHIC20n1 => return "L4PHIC20n1";
       when L4PHID32n2 => return "L4PHID32n2";
       when L4PHIB9n1 => return "L4PHIB9n1";
       when L4PHIA7n3 => return "L4PHIA7n3";
       when L6PHIB14n1 => return "L6PHIB14n1";
       when L4PHID30n2 => return "L4PHID30n2";
       when L4PHIA4n2 => return "L4PHIA4n2";
       when L6PHIA6n1 => return "L6PHIA6n1";
       when L4PHID29n1 => return "L4PHID29n1";
       when L4PHIA6n3 => return "L4PHIA6n3";
       when L6PHID31n1 => return "L6PHID31n1";
       when L6PHIA4n3 => return "L6PHIA4n3";
       when L6PHIC18n4 => return "L6PHIC18n4";
       when L6PHID29n3 => return "L6PHID29n3";
       when L6PHIC17n2 => return "L6PHIC17n2";
       when L4PHID27n3 => return "L4PHID27n3";
       when L4PHIC20n3 => return "L4PHIC20n3";
       when L4PHIC19n2 => return "L4PHIC19n2";
       when L4PHIB10n3 => return "L4PHIB10n3";
       when L4PHIC19n3 => return "L4PHIC19n3";
       when L6PHIA1n2 => return "L6PHIA1n2";
       when L6PHIA7n2 => return "L6PHIA7n2";
       when L6PHIC23n1 => return "L6PHIC23n1";
       when L4PHIB15n3 => return "L4PHIB15n3";
       when L6PHIB16n2 => return "L6PHIB16n2";
       when L6PHIC20n1 => return "L6PHIC20n1";
       when L4PHIC17n2 => return "L4PHIC17n2";
       when L4PHIB12n3 => return "L4PHIB12n3";
       when L6PHIA8n4 => return "L6PHIA8n4";
       when L6PHIC23n2 => return "L6PHIC23n2";
       when L4PHIC21n3 => return "L4PHIC21n3";
       when L4PHIB10n1 => return "L4PHIB10n1";
       when L6PHIA7n1 => return "L6PHIA7n1";
       when L6PHIC20n3 => return "L6PHIC20n3";
       when L4PHIB15n1 => return "L4PHIB15n1";
       when L6PHID26n3 => return "L6PHID26n3";
       when L6PHIC22n2 => return "L6PHIC22n2";
       when L4PHID28n3 => return "L4PHID28n3";
       when L6PHIA5n1 => return "L6PHIA5n1";
       when L6PHID32n1 => return "L6PHID32n1";
       when L4PHID26n3 => return "L4PHID26n3";
       when L6PHIB11n2 => return "L6PHIB11n2";
       when L6PHIA4n1 => return "L6PHIA4n1";
       when L4PHID30n3 => return "L4PHID30n3";
       when L4PHID29n2 => return "L4PHID29n2";
       when L6PHIC23n3 => return "L6PHIC23n3";
       when L6PHIC18n3 => return "L6PHIC18n3";
       when L6PHIA8n2 => return "L6PHIA8n2";
       when L6PHIA3n2 => return "L6PHIA3n2";
       when L4PHID26n2 => return "L4PHID26n2";
       when L4PHID28n2 => return "L4PHID28n2";
       when L4PHID31n2 => return "L4PHID31n2";
       when L6PHIB16n1 => return "L6PHIB16n1";
       when L6PHID31n3 => return "L6PHID31n3";
       when L6PHIC18n2 => return "L6PHIC18n2";
       when L4PHIB9n2 => return "L4PHIB9n2";
       when L4PHIA8n1 => return "L4PHIA8n1";
       when L4PHIC23n1 => return "L4PHIC23n1";
       when L6PHID27n3 => return "L6PHID27n3";
       when L4PHID32n1 => return "L4PHID32n1";
       when L4PHIB11n1 => return "L4PHIB11n1";
       when L6PHID26n4 => return "L6PHID26n4";
       when L6PHID31n2 => return "L6PHID31n2";
       when L6PHIA2n2 => return "L6PHIA2n2";
       when L6PHIC21n3 => return "L6PHIC21n3";
       when L4PHIB12n1 => return "L4PHIB12n1";
       when L6PHID32n2 => return "L6PHID32n2";
       when L6PHID25n4 => return "L6PHID25n4";
       when L6PHIA2n1 => return "L6PHIA2n1";
       when L4PHIA5n3 => return "L4PHIA5n3";
       when L6PHID28n4 => return "L6PHID28n4";
       when L4PHIC23n2 => return "L4PHIC23n2";
       when L4PHIB12n2 => return "L4PHIB12n2";
       when L6PHIB10n1 => return "L6PHIB10n1";
       when L4PHIC21n2 => return "L4PHIC21n2";
       when L6PHIB10n2 => return "L6PHIB10n2";
       when L4PHIC24n1 => return "L4PHIC24n1";
       when L6PHIA6n2 => return "L6PHIA6n2";
       when L6PHIC22n3 => return "L6PHIC22n3";
       when L6PHIB13n1 => return "L6PHIB13n1";
       when L4PHIB9n3 => return "L4PHIB9n3";
       when L4PHIB16n1 => return "L4PHIB16n1";
       when L6PHID30n1 => return "L6PHID30n1";
       when L4PHID29n3 => return "L4PHID29n3";
       when L6PHIA6n4 => return "L6PHIA6n4";
       when L6PHIB15n2 => return "L6PHIB15n2";
       when L4PHID30n1 => return "L4PHID30n1";
       when L6PHIC20n4 => return "L6PHIC20n4";
       when L6PHIC22n4 => return "L6PHIC22n4";
       when L6PHIB15n4 => return "L6PHIB15n4";
       when L4PHIB16n3 => return "L4PHIB16n3";
       when L4PHIC19n1 => return "L4PHIC19n1";
       when L4PHIA2n1 => return "L4PHIA2n1";
       when L6PHIC19n4 => return "L6PHIC19n4";
       when L6PHIC21n2 => return "L6PHIC21n2";
       when L6PHIC21n1 => return "L6PHIC21n1";
       when L4PHIB14n1 => return "L4PHIB14n1";
       when L6PHIB16n4 => return "L6PHIB16n4";
       when L4PHIA6n2 => return "L4PHIA6n2";
       when L4PHID26n1 => return "L4PHID26n1";
       when L6PHIC24n1 => return "L6PHIC24n1";
       when L4PHIA8n2 => return "L4PHIA8n2";
       when L6PHIA3n1 => return "L6PHIA3n1";
       when L6PHIA4n4 => return "L6PHIA4n4";
       when L6PHIB9n3 => return "L6PHIB9n3";
       when L6PHIB10n4 => return "L6PHIB10n4";
       when L4PHIB13n1 => return "L4PHIB13n1";
       when L4PHID25n3 => return "L4PHID25n3";
       when L6PHIA2n3 => return "L6PHIA2n3";
       when L6PHID29n2 => return "L6PHID29n2";
       when L4PHIC22n1 => return "L4PHIC22n1";
       when L6PHIC20n2 => return "L6PHIC20n2";
       when L4PHIC23n3 => return "L4PHIC23n3";
       when L6PHIC23n4 => return "L6PHIC23n4";
       when L4PHIA3n3 => return "L4PHIA3n3";
       when L4PHIC17n1 => return "L4PHIC17n1";
       when L6PHIB13n3 => return "L6PHIB13n3";
       when L4PHIA4n3 => return "L4PHIA4n3";
       when L4PHIA3n1 => return "L4PHIA3n1";
       when L6PHID30n2 => return "L6PHID30n2";
       when L4PHIA8n3 => return "L4PHIA8n3";
       when L4PHIA7n2 => return "L4PHIA7n2";
       when L6PHIC17n1 => return "L6PHIC17n1";
       when L4PHIA1n1 => return "L4PHIA1n1";
       when L4PHID27n2 => return "L4PHID27n2";
       when L4PHIA1n2 => return "L4PHIA1n2";
       when L6PHIA5n3 => return "L6PHIA5n3";
       when L6PHID26n2 => return "L6PHID26n2";
       when L6PHIC24n3 => return "L6PHIC24n3";
       when L4PHIA2n2 => return "L4PHIA2n2";
       when L6PHID30n3 => return "L6PHID30n3";
       when L4PHIC24n3 => return "L4PHIC24n3";
       when L4PHID28n1 => return "L4PHID28n1";
       when L6PHIB14n4 => return "L6PHIB14n4";
       when L6PHIB9n1 => return "L6PHIB9n1";
       when L6PHIC24n4 => return "L6PHIC24n4";
       when L6PHIA1n1 => return "L6PHIA1n1";
       when L4PHIB15n2 => return "L4PHIB15n2";
       when L6PHIB16n3 => return "L6PHIB16n3";
       when L6PHIA5n4 => return "L6PHIA5n4";
       when L4PHID31n1 => return "L4PHID31n1";
       when L4PHIA5n2 => return "L4PHIA5n2";
       when L6PHIA5n2 => return "L6PHIA5n2";
       when L6PHIB13n4 => return "L6PHIB13n4";
       when L4PHIB11n2 => return "L4PHIB11n2";
       when L4PHID27n1 => return "L4PHID27n1";
       when L4PHIA3n2 => return "L4PHIA3n2";
       when L4PHIC21n1 => return "L4PHIC21n1";
       when L6PHIA4n2 => return "L6PHIA4n2";
       when L4PHIA7n1 => return "L4PHIA7n1";
       when L6PHIC17n4 => return "L6PHIC17n4";
       when L4PHIC18n2 => return "L4PHIC18n2";
       when L4PHIB11n3 => return "L4PHIB11n3";
       when L6PHIB12n3 => return "L6PHIB12n3";
       when L6PHIC21n4 => return "L6PHIC21n4";
       when L4PHIC24n2 => return "L4PHIC24n2";
       when L4PHIA5n1 => return "L4PHIA5n1";
       when L6PHIB9n4 => return "L6PHIB9n4";
       when L4PHIB10n2 => return "L4PHIB10n2";
       when L4PHIC22n3 => return "L4PHIC22n3";
       when L6PHIA8n1 => return "L6PHIA8n1";
       when L6PHID28n3 => return "L6PHID28n3";
       when L6PHIC19n3 => return "L6PHIC19n3";
       when L6PHIA7n4 => return "L6PHIA7n4";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSTE_23) return string is
  begin
    case val is
       when L5PHIB7n1 => return "L5PHIB7n1";
       when L5PHIC10n3 => return "L5PHIC10n3";
       when L5PHID15n1 => return "L5PHID15n1";
       when L5PHIB6n4 => return "L5PHIB6n4";
       when L5PHIB8n8 => return "L5PHIB8n8";
       when L5PHIC12n6 => return "L5PHIC12n6";
       when L5PHID16n5 => return "L5PHID16n5";
       when L5PHIC11n5 => return "L5PHIC11n5";
       when L5PHID15n3 => return "L5PHID15n3";
       when L5PHIA3n7 => return "L5PHIA3n7";
       when L5PHID14n2 => return "L5PHID14n2";
       when L5PHID13n5 => return "L5PHID13n5";
       when L5PHIA4n8 => return "L5PHIA4n8";
       when L5PHIB8n7 => return "L5PHIB8n7";
       when L5PHIA3n5 => return "L5PHIA3n5";
       when L5PHIB5n3 => return "L5PHIB5n3";
       when L5PHIC12n2 => return "L5PHIC12n2";
       when L5PHIB8n4 => return "L5PHIB8n4";
       when L5PHIC9n1 => return "L5PHIC9n1";
       when L5PHIC10n8 => return "L5PHIC10n8";
       when L5PHID16n2 => return "L5PHID16n2";
       when L5PHIC12n5 => return "L5PHIC12n5";
       when L5PHIB6n2 => return "L5PHIB6n2";
       when L5PHIC9n4 => return "L5PHIC9n4";
       when L5PHIA1n1 => return "L5PHIA1n1";
       when L5PHIB7n8 => return "L5PHIB7n8";
       when L5PHIA4n4 => return "L5PHIA4n4";
       when L5PHIB7n4 => return "L5PHIB7n4";
       when L5PHID13n3 => return "L5PHID13n3";
       when L5PHIB6n1 => return "L5PHIB6n1";
       when L5PHID15n4 => return "L5PHID15n4";
       when L5PHIC11n1 => return "L5PHIC11n1";
       when L5PHIA4n6 => return "L5PHIA4n6";
       when L5PHIC12n4 => return "L5PHIC12n4";
       when L5PHIC11n2 => return "L5PHIC11n2";
       when L5PHIA3n4 => return "L5PHIA3n4";
       when L5PHID13n4 => return "L5PHID13n4";
       when L5PHID13n2 => return "L5PHID13n2";
       when L5PHIB5n8 => return "L5PHIB5n8";
       when L5PHIC9n3 => return "L5PHIC9n3";
       when L5PHIA3n6 => return "L5PHIA3n6";
       when L5PHID14n5 => return "L5PHID14n5";
       when L5PHIC11n8 => return "L5PHIC11n8";
       when L5PHIA2n6 => return "L5PHIA2n6";
       when L5PHIB8n3 => return "L5PHIB8n3";
       when L5PHIC11n4 => return "L5PHIC11n4";
       when L5PHIC12n1 => return "L5PHIC12n1";
       when L5PHIA1n2 => return "L5PHIA1n2";
       when L5PHIB7n2 => return "L5PHIB7n2";
       when L5PHIA2n7 => return "L5PHIA2n7";
       when L5PHIA3n2 => return "L5PHIA3n2";
       when L5PHIA4n2 => return "L5PHIA4n2";
       when L5PHIB5n2 => return "L5PHIB5n2";
       when L5PHIA3n8 => return "L5PHIA3n8";
       when L5PHIC11n6 => return "L5PHIC11n6";
       when L5PHID14n4 => return "L5PHID14n4";
       when L5PHIA2n2 => return "L5PHIA2n2";
       when L5PHID16n1 => return "L5PHID16n1";
       when L5PHID13n7 => return "L5PHID13n7";
       when L5PHIA2n5 => return "L5PHIA2n5";
       when L5PHID14n7 => return "L5PHID14n7";
       when L5PHIC12n8 => return "L5PHIC12n8";
       when L5PHIA2n4 => return "L5PHIA2n4";
       when L5PHID13n1 => return "L5PHID13n1";
       when L5PHIB7n5 => return "L5PHIB7n5";
       when L5PHIC10n7 => return "L5PHIC10n7";
       when L5PHIA1n4 => return "L5PHIA1n4";
       when L5PHIC9n6 => return "L5PHIC9n6";
       when L5PHID16n4 => return "L5PHID16n4";
       when L5PHIA2n1 => return "L5PHIA2n1";
       when L5PHIC10n2 => return "L5PHIC10n2";
       when L5PHIA4n3 => return "L5PHIA4n3";
       when L5PHIC12n3 => return "L5PHIC12n3";
       when L5PHIB7n3 => return "L5PHIB7n3";
       when L5PHIB6n8 => return "L5PHIB6n8";
       when L5PHIB8n1 => return "L5PHIB8n1";
       when L5PHIB6n3 => return "L5PHIB6n3";
       when L5PHIA2n3 => return "L5PHIA2n3";
       when L5PHIC12n7 => return "L5PHIC12n7";
       when L5PHIC11n7 => return "L5PHIC11n7";
       when L5PHIC9n5 => return "L5PHIC9n5";
       when L5PHIC9n7 => return "L5PHIC9n7";
       when L5PHID13n8 => return "L5PHID13n8";
       when L5PHIC11n3 => return "L5PHIC11n3";
       when L5PHIC9n2 => return "L5PHIC9n2";
       when L5PHIC10n1 => return "L5PHIC10n1";
       when L5PHIB5n6 => return "L5PHIB5n6";
       when L5PHIC10n5 => return "L5PHIC10n5";
       when L5PHIB5n1 => return "L5PHIB5n1";
       when L5PHIA3n1 => return "L5PHIA3n1";
       when L5PHIA4n7 => return "L5PHIA4n7";
       when L5PHID14n3 => return "L5PHID14n3";
       when L5PHIC10n4 => return "L5PHIC10n4";
       when L5PHIB8n2 => return "L5PHIB8n2";
       when L5PHIA1n5 => return "L5PHIA1n5";
       when L5PHIB5n5 => return "L5PHIB5n5";
       when L5PHID15n7 => return "L5PHID15n7";
       when L5PHIA3n3 => return "L5PHIA3n3";
       when L5PHID16n3 => return "L5PHID16n3";
       when L5PHID14n1 => return "L5PHID14n1";
       when L5PHIB5n7 => return "L5PHIB5n7";
       when L5PHIB6n6 => return "L5PHIB6n6";
       when L5PHIA4n1 => return "L5PHIA4n1";
       when L5PHIB8n6 => return "L5PHIB8n6";
       when L5PHID14n6 => return "L5PHID14n6";
       when L5PHID15n2 => return "L5PHID15n2";
       when L5PHIA4n5 => return "L5PHIA4n5";
       when L5PHIB6n5 => return "L5PHIB6n5";
       when L5PHID15n6 => return "L5PHID15n6";
       when L5PHIB7n7 => return "L5PHIB7n7";
       when L5PHID15n5 => return "L5PHID15n5";
       when L5PHIC9n8 => return "L5PHIC9n8";
       when L5PHID14n8 => return "L5PHID14n8";
       when L5PHID13n6 => return "L5PHID13n6";
       when L5PHIB7n6 => return "L5PHIB7n6";
       when L5PHIC10n6 => return "L5PHIC10n6";
       when L5PHIB8n5 => return "L5PHIB8n5";
       when L5PHIA1n3 => return "L5PHIA1n3";
       when L5PHIB5n4 => return "L5PHIB5n4";
       when L5PHIB6n7 => return "L5PHIB6n7";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMSTE_16) return string is
  begin
    case val is
       when L2PHID28n3 => return "L2PHID28n3";
       when L2PHID30n1 => return "L2PHID30n1";
       when L2PHID27n2 => return "L2PHID27n2";
       when L2PHIC23n3 => return "L2PHIC23n3";
       when L2PHIB13n3 => return "L2PHIB13n3";
       when L3PHIJ7n3 => return "L3PHIJ7n3";
       when L2PHIA8n4 => return "L2PHIA8n4";
       when L3PHIJ8n1 => return "L3PHIJ8n1";
       when L2PHIB9n5 => return "L2PHIB9n5";
       when L2PHIC20n5 => return "L2PHIC20n5";
       when L2PHIC22n1 => return "L2PHIC22n1";
       when L2PHIB10n1 => return "L2PHIB10n1";
       when L3PHII1n1 => return "L3PHII1n1";
       when L2PHIB12n3 => return "L2PHIB12n3";
       when L2PHIB9n4 => return "L2PHIB9n4";
       when L3PHIK9n3 => return "L3PHIK9n3";
       when L2PHIC22n2 => return "L2PHIC22n2";
       when L2PHID32n2 => return "L2PHID32n2";
       when L2PHIC24n1 => return "L2PHIC24n1";
       when L2PHID30n4 => return "L2PHID30n4";
       when L3PHII3n3 => return "L3PHII3n3";
       when L3PHII1n2 => return "L3PHII1n2";
       when L2PHID30n2 => return "L2PHID30n2";
       when L3PHIK11n2 => return "L3PHIK11n2";
       when L2PHIC22n4 => return "L2PHIC22n4";
       when L2PHIA2n2 => return "L2PHIA2n2";
       when L3PHIL14n3 => return "L3PHIL14n3";
       when L2PHIB16n3 => return "L2PHIB16n3";
       when L2PHID30n3 => return "L2PHID30n3";
       when L2PHIA4n2 => return "L2PHIA4n2";
       when L2PHID28n2 => return "L2PHID28n2";
       when L3PHIK10n2 => return "L3PHIK10n2";
       when L2PHIC18n1 => return "L2PHIC18n1";
       when L2PHIB15n1 => return "L2PHIB15n1";
       when L2PHIC22n3 => return "L2PHIC22n3";
       when L2PHIC22n5 => return "L2PHIC22n5";
       when L2PHID32n3 => return "L2PHID32n3";
       when L2PHIB14n4 => return "L2PHIB14n4";
       when L2PHIA4n3 => return "L2PHIA4n3";
       when L2PHIB16n2 => return "L2PHIB16n2";
       when L3PHIJ8n3 => return "L3PHIJ8n3";
       when L2PHIB16n4 => return "L2PHIB16n4";
       when L2PHIB15n4 => return "L2PHIB15n4";
       when L2PHIA3n3 => return "L2PHIA3n3";
       when L2PHIB10n2 => return "L2PHIB10n2";
       when L3PHIJ5n3 => return "L3PHIJ5n3";
       when L2PHIB12n1 => return "L2PHIB12n1";
       when L2PHIC21n2 => return "L2PHIC21n2";
       when L2PHID27n3 => return "L2PHID27n3";
       when L2PHIA5n1 => return "L2PHIA5n1";
       when L2PHIB12n5 => return "L2PHIB12n5";
       when L2PHID25n2 => return "L2PHID25n2";
       when L2PHIC23n5 => return "L2PHIC23n5";
       when L2PHIB11n3 => return "L2PHIB11n3";
       when L3PHIJ6n3 => return "L3PHIJ6n3";
       when L2PHIC17n4 => return "L2PHIC17n4";
       when L2PHIB10n5 => return "L2PHIB10n5";
       when L3PHIL15n1 => return "L3PHIL15n1";
       when L2PHIA8n3 => return "L2PHIA8n3";
       when L3PHIK9n2 => return "L3PHIK9n2";
       when L3PHII4n3 => return "L3PHII4n3";
       when L2PHIA4n1 => return "L2PHIA4n1";
       when L2PHIA7n5 => return "L2PHIA7n5";
       when L2PHID27n4 => return "L2PHID27n4";
       when L2PHIA1n1 => return "L2PHIA1n1";
       when L2PHID29n1 => return "L2PHID29n1";
       when L2PHIC23n1 => return "L2PHIC23n1";
       when L2PHIA2n1 => return "L2PHIA2n1";
       when L2PHIC19n2 => return "L2PHIC19n2";
       when L2PHID29n2 => return "L2PHID29n2";
       when L2PHIC23n4 => return "L2PHIC23n4";
       when L2PHID26n3 => return "L2PHID26n3";
       when L2PHIA3n1 => return "L2PHIA3n1";
       when L2PHIB11n4 => return "L2PHIB11n4";
       when L2PHIC18n5 => return "L2PHIC18n5";
       when L3PHIL15n3 => return "L3PHIL15n3";
       when L2PHID25n3 => return "L2PHID25n3";
       when L2PHIC17n1 => return "L2PHIC17n1";
       when L2PHID28n4 => return "L2PHID28n4";
       when L2PHIC17n2 => return "L2PHIC17n2";
       when L2PHIC24n5 => return "L2PHIC24n5";
       when L2PHIC19n1 => return "L2PHIC19n1";
       when L2PHIB12n4 => return "L2PHIB12n4";
       when L2PHIC24n3 => return "L2PHIC24n3";
       when L3PHII2n1 => return "L3PHII2n1";
       when L2PHIA1n2 => return "L2PHIA1n2";
       when L2PHID28n1 => return "L2PHID28n1";
       when L2PHIB13n2 => return "L2PHIB13n2";
       when L2PHID26n1 => return "L2PHID26n1";
       when L2PHIC20n2 => return "L2PHIC20n2";
       when L3PHIL13n2 => return "L3PHIL13n2";
       when L2PHID26n5 => return "L2PHID26n5";
       when L2PHIA5n3 => return "L2PHIA5n3";
       when L2PHIB10n4 => return "L2PHIB10n4";
       when L2PHIA8n5 => return "L2PHIA8n5";
       when L3PHIJ7n1 => return "L3PHIJ7n1";
       when L2PHIA7n4 => return "L2PHIA7n4";
       when L2PHID27n5 => return "L2PHID27n5";
       when L3PHII3n1 => return "L3PHII3n1";
       when L2PHIC18n2 => return "L2PHIC18n2";
       when L2PHIA3n2 => return "L2PHIA3n2";
       when L3PHIK11n3 => return "L3PHIK11n3";
       when L2PHIA5n4 => return "L2PHIA5n4";
       when L2PHIA4n4 => return "L2PHIA4n4";
       when L2PHIC21n3 => return "L2PHIC21n3";
       when L2PHIA2n4 => return "L2PHIA2n4";
       when L3PHIK10n3 => return "L3PHIK10n3";
       when L2PHIC19n4 => return "L2PHIC19n4";
       when L2PHIB11n1 => return "L2PHIB11n1";
       when L2PHIA6n3 => return "L2PHIA6n3";
       when L2PHIB14n5 => return "L2PHIB14n5";
       when L2PHIB9n1 => return "L2PHIB9n1";
       when L3PHIK12n3 => return "L3PHIK12n3";
       when L2PHIB15n3 => return "L2PHIB15n3";
       when L2PHID32n1 => return "L2PHID32n1";
       when L2PHIC19n3 => return "L2PHIC19n3";
       when L3PHIJ8n2 => return "L3PHIJ8n2";
       when L3PHIK12n2 => return "L3PHIK12n2";
       when L2PHIA5n5 => return "L2PHIA5n5";
       when L2PHIA1n3 => return "L2PHIA1n3";
       when L2PHIB14n2 => return "L2PHIB14n2";
       when L2PHIC21n5 => return "L2PHIC21n5";
       when L3PHIL15n2 => return "L3PHIL15n2";
       when L2PHID26n2 => return "L2PHID26n2";
       when L2PHIA6n2 => return "L2PHIA6n2";
       when L3PHII3n2 => return "L3PHII3n2";
       when L2PHIB10n3 => return "L2PHIB10n3";
       when L2PHIB13n5 => return "L2PHIB13n5";
       when L3PHII2n2 => return "L3PHII2n2";
       when L3PHIJ7n2 => return "L3PHIJ7n2";
       when L2PHIC20n3 => return "L2PHIC20n3";
       when L3PHII4n1 => return "L3PHII4n1";
       when L2PHID26n4 => return "L2PHID26n4";
       when L2PHIA7n1 => return "L2PHIA7n1";
       when L2PHIA8n2 => return "L2PHIA8n2";
       when L2PHIB11n2 => return "L2PHIB11n2";
       when L2PHIC21n1 => return "L2PHIC21n1";
       when L2PHID31n3 => return "L2PHID31n3";
       when L2PHIC17n3 => return "L2PHIC17n3";
       when L2PHID27n1 => return "L2PHID27n1";
       when L2PHID29n5 => return "L2PHID29n5";
       when L2PHID31n2 => return "L2PHID31n2";
       when L2PHIB9n3 => return "L2PHIB9n3";
       when L2PHIB15n2 => return "L2PHIB15n2";
       when L2PHIC18n3 => return "L2PHIC18n3";
       when L3PHIL13n3 => return "L3PHIL13n3";
       when L2PHIA7n2 => return "L2PHIA7n2";
       when L2PHIA3n4 => return "L2PHIA3n4";
       when L2PHID31n4 => return "L2PHID31n4";
       when L2PHIC20n4 => return "L2PHIC20n4";
       when L2PHIC19n5 => return "L2PHIC19n5";
       when L2PHIB13n1 => return "L2PHIB13n1";
       when L2PHIB12n2 => return "L2PHIB12n2";
       when L2PHIB13n4 => return "L2PHIB13n4";
       when L3PHIL16n2 => return "L3PHIL16n2";
       when L3PHIL14n2 => return "L3PHIL14n2";
       when L2PHIA5n2 => return "L2PHIA5n2";
       when L3PHIJ6n2 => return "L3PHIJ6n2";
       when L2PHIC24n4 => return "L2PHIC24n4";
       when L2PHIA6n5 => return "L2PHIA6n5";
       when L2PHIC17n5 => return "L2PHIC17n5";
       when L3PHIL13n1 => return "L3PHIL13n1";
       when L3PHIL16n1 => return "L3PHIL16n1";
       when L2PHIA8n1 => return "L2PHIA8n1";
       when L2PHID25n1 => return "L2PHID25n1";
       when L2PHIA4n5 => return "L2PHIA4n5";
       when L2PHIB16n5 => return "L2PHIB16n5";
       when L2PHIB14n3 => return "L2PHIB14n3";
       when L2PHID28n5 => return "L2PHID28n5";
       when L2PHID25n5 => return "L2PHID25n5";
       when L2PHID29n4 => return "L2PHID29n4";
       when L2PHIB14n1 => return "L2PHIB14n1";
       when L2PHIA2n3 => return "L2PHIA2n3";
       when L3PHII4n2 => return "L3PHII4n2";
       when L2PHIB11n5 => return "L2PHIB11n5";
       when L2PHIB15n5 => return "L2PHIB15n5";
       when L2PHIA7n3 => return "L2PHIA7n3";
       when L2PHIC18n4 => return "L2PHIC18n4";
       when L3PHIL14n1 => return "L3PHIL14n1";
       when L2PHID29n3 => return "L2PHID29n3";
       when L2PHID30n5 => return "L2PHID30n5";
       when L3PHIK10n1 => return "L3PHIK10n1";
       when L3PHIK11n1 => return "L3PHIK11n1";
       when L2PHIA6n4 => return "L2PHIA6n4";
       when L2PHID31n1 => return "L2PHID31n1";
       when L3PHIJ5n1 => return "L3PHIJ5n1";
       when L2PHIA6n1 => return "L2PHIA6n1";
       when L2PHIC20n1 => return "L2PHIC20n1";
       when L2PHIC23n2 => return "L2PHIC23n2";
       when L3PHIJ5n2 => return "L3PHIJ5n2";
       when L2PHIC24n2 => return "L2PHIC24n2";
       when L3PHIJ6n1 => return "L3PHIJ6n1";
       when L2PHIB16n1 => return "L2PHIB16n1";
       when L2PHIB9n2 => return "L2PHIB9n2";
       when L2PHID25n4 => return "L2PHID25n4";
       when L2PHIA3n5 => return "L2PHIA3n5";
       when L3PHIK9n1 => return "L3PHIK9n1";
       when L2PHIC21n4 => return "L2PHIC21n4";
       when L3PHII2n3 => return "L3PHII2n3";
       when L3PHIK12n1 => return "L3PHIK12n1";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_SP_14) return string is
  begin
    case val is
       when L3PHID14_L4PHID29 => return "L3PHID14_L4PHID29";
       when L3PHID14_L4PHID25 => return "L3PHID14_L4PHID25";
       when L1PHIF21_L2PHIC22 => return "L1PHIF21_L2PHIC22";
       when L1PHIE18_L2PHIB16 => return "L1PHIE18_L2PHIB16";
       when L3PHIC9_L4PHIC17 => return "L3PHIC9_L4PHIC17";
       when L5PHIA1_L6PHIA2 => return "L5PHIA1_L6PHIA2";
       when L3PHID13_L4PHID26 => return "L3PHID13_L4PHID26";
       when L2PHII4_L3PHII4 => return "L2PHII4_L3PHII4";
       when L5PHIC11_L6PHIC23 => return "L5PHIC11_L6PHIC23";
       when L2PHIK12_L3PHIK12 => return "L2PHIK12_L3PHIK12";
       when L5PHIB6_L6PHIB10 => return "L5PHIB6_L6PHIB10";
       when L3PHIA1_L4PHIA3 => return "L3PHIA1_L4PHIA3";
       when L3PHIA1_L4PHIA1 => return "L3PHIA1_L4PHIA1";
       when L1PHIA2_L2PHIA2 => return "L1PHIA2_L2PHIA2";
       when L3PHIB5_L4PHIA8 => return "L3PHIB5_L4PHIA8";
       when L3PHIC11_L4PHIC20 => return "L3PHIC11_L4PHIC20";
       when L1PHIG26_L2PHID27 => return "L1PHIG26_L2PHID27";
       when L5PHID14_L6PHID26 => return "L5PHID14_L6PHID26";
       when L1PHIH31_L2PHID29 => return "L1PHIH31_L2PHID29";
       when L1PHIC10_L2PHIB9 => return "L1PHIC10_L2PHIB9";
       when L1PHIC12_L2PHIB12 => return "L1PHIC12_L2PHIB12";
       when L3PHIB8_L4PHIB14 => return "L3PHIB8_L4PHIB14";
       when L3PHIA3_L4PHIA5 => return "L3PHIA3_L4PHIA5";
       when L1PHIF23_L2PHID25 => return "L1PHIF23_L2PHID25";
       when L2PHIJ5_L3PHIJ5 => return "L2PHIJ5_L3PHIJ5";
       when L5PHIA3_L6PHIA6 => return "L5PHIA3_L6PHIA6";
       when L1PHIE19_L2PHIC17 => return "L1PHIE19_L2PHIC17";
       when L3PHIB7_L4PHIB11 => return "L3PHIB7_L4PHIB11";
       when L2PHII3_L3PHII3 => return "L2PHII3_L3PHII3";
       when L5PHIB8_L6PHIC18 => return "L5PHIB8_L6PHIC18";
       when L1PHIG25_L2PHID26 => return "L1PHIG25_L2PHID26";
       when L1PHIB7_L2PHIB9 => return "L1PHIB7_L2PHIB9";
       when L1PHIA4_L2PHIA6 => return "L1PHIA4_L2PHIA6";
       when L3PHIA4_L4PHIA5 => return "L3PHIA4_L4PHIA5";
       when L1PHIE17_L2PHIB16 => return "L1PHIE17_L2PHIB16";
       when L1PHID15_L2PHIC17 => return "L1PHID15_L2PHIC17";
       when L5PHID13_L6PHID27 => return "L5PHID13_L6PHID27";
       when L5PHIB8_L6PHIB13 => return "L5PHIB8_L6PHIB13";
       when L1PHIF24_L2PHIC24 => return "L1PHIF24_L2PHIC24";
       when L1PHIG26_L2PHID28 => return "L1PHIG26_L2PHID28";
       when L3PHIC11_L4PHIC24 => return "L3PHIC11_L4PHIC24";
       when L2PHII3_L3PHII2 => return "L2PHII3_L3PHII2";
       when L1PHIG28_L2PHID30 => return "L1PHIG28_L2PHID30";
       when L5PHIB8_L6PHIB14 => return "L5PHIB8_L6PHIB14";
       when L5PHIB6_L6PHIB13 => return "L5PHIB6_L6PHIB13";
       when L3PHIA3_L4PHIA3 => return "L3PHIA3_L4PHIA3";
       when L1PHIF21_L2PHIC21 => return "L1PHIF21_L2PHIC21";
       when L2PHIK10_L3PHIK10 => return "L2PHIK10_L3PHIK10";
       when L5PHIB5_L6PHIB12 => return "L5PHIB5_L6PHIB12";
       when L5PHIC12_L6PHIC21 => return "L5PHIC12_L6PHIC21";
       when L3PHIA3_L4PHIA4 => return "L3PHIA3_L4PHIA4";
       when L5PHIC12_L6PHIC24 => return "L5PHIC12_L6PHIC24";
       when L3PHIC12_L4PHIC22 => return "L3PHIC12_L4PHIC22";
       when L1PHIA1_L2PHIA3 => return "L1PHIA1_L2PHIA3";
       when L5PHID16_L6PHID29 => return "L5PHID16_L6PHID29";
       when L5PHID16_L6PHID32 => return "L5PHID16_L6PHID32";
       when L3PHIC12_L4PHIC21 => return "L3PHIC12_L4PHIC21";
       when L5PHID15_L6PHID29 => return "L5PHID15_L6PHID29";
       when L3PHIA4_L4PHIA8 => return "L3PHIA4_L4PHIA8";
       when L3PHIB5_L4PHIA7 => return "L3PHIB5_L4PHIA7";
       when L5PHID14_L6PHID28 => return "L5PHID14_L6PHID28";
       when L2PHIL15_L3PHIL14 => return "L2PHIL15_L3PHIL14";
       when L5PHIC12_L6PHIC23 => return "L5PHIC12_L6PHIC23";
       when L3PHIA1_L4PHIA4 => return "L3PHIA1_L4PHIA4";
       when L1PHID16_L2PHIB15 => return "L1PHID16_L2PHIB15";
       when L1PHIC10_L2PHIB11 => return "L1PHIC10_L2PHIB11";
       when L1PHIF24_L2PHIC22 => return "L1PHIF24_L2PHIC22";
       when L3PHIA3_L4PHIA7 => return "L3PHIA3_L4PHIA7";
       when L5PHIA4_L6PHIA6 => return "L5PHIA4_L6PHIA6";
       when L5PHID13_L6PHID29 => return "L5PHID13_L6PHID29";
       when L5PHIC12_L6PHIC20 => return "L5PHIC12_L6PHIC20";
       when L3PHIA2_L4PHIA2 => return "L3PHIA2_L4PHIA2";
       when L1PHIH30_L2PHID30 => return "L1PHIH30_L2PHID30";
       when L5PHIC10_L6PHIC18 => return "L5PHIC10_L6PHIC18";
       when L5PHIC11_L6PHIC18 => return "L5PHIC11_L6PHIC18";
       when L1PHIE18_L2PHIC20 => return "L1PHIE18_L2PHIC20";
       when L3PHIC11_L4PHIC21 => return "L3PHIC11_L4PHIC21";
       when L3PHIA4_L4PHIA7 => return "L3PHIA4_L4PHIA7";
       when L3PHID13_L4PHID25 => return "L3PHID13_L4PHID25";
       when L3PHIC12_L4PHIC23 => return "L3PHIC12_L4PHIC23";
       when L1PHIC9_L2PHIB9 => return "L1PHIC9_L2PHIB9";
       when L5PHIA4_L6PHIA8 => return "L5PHIA4_L6PHIA8";
       when L1PHIA4_L2PHIA5 => return "L1PHIA4_L2PHIA5";
       when L1PHID16_L2PHIB14 => return "L1PHID16_L2PHIB14";
       when L3PHIB6_L4PHIB10 => return "L3PHIB6_L4PHIB10";
       when L5PHID14_L6PHID31 => return "L5PHID14_L6PHID31";
       when L1PHIH32_L2PHID32 => return "L1PHIH32_L2PHID32";
       when L2PHIL14_L3PHIL15 => return "L2PHIL14_L3PHIL15";
       when L3PHIA2_L4PHIA1 => return "L3PHIA2_L4PHIA1";
       when L2PHIK12_L3PHIL13 => return "L2PHIK12_L3PHIL13";
       when L3PHIC9_L4PHIC19 => return "L3PHIC9_L4PHIC19";
       when L3PHIA4_L4PHIA6 => return "L3PHIA4_L4PHIA6";
       when L5PHIC12_L6PHID27 => return "L5PHIC12_L6PHID27";
       when L1PHIE19_L2PHIC20 => return "L1PHIE19_L2PHIC20";
       when L3PHIC10_L4PHIC21 => return "L3PHIC10_L4PHIC21";
       when L1PHIB8_L2PHIB10 => return "L1PHIB8_L2PHIB10";
       when L1PHIG28_L2PHID29 => return "L1PHIG28_L2PHID29";
       when L1PHIB5_L2PHIA6 => return "L1PHIB5_L2PHIA6";
       when L5PHIC10_L6PHIC20 => return "L5PHIC10_L6PHIC20";
       when L1PHIA3_L2PHIA2 => return "L1PHIA3_L2PHIA2";
       when L5PHIB6_L6PHIB12 => return "L5PHIB6_L6PHIB12";
       when L5PHIB8_L6PHIC19 => return "L5PHIB8_L6PHIC19";
       when L2PHII1_L3PHII2 => return "L2PHII1_L3PHII2";
       when L5PHIB8_L6PHIB12 => return "L5PHIB8_L6PHIB12";
       when L5PHIA3_L6PHIA5 => return "L5PHIA3_L6PHIA5";
       when L1PHIG27_L2PHID28 => return "L1PHIG27_L2PHID28";
       when L1PHIC12_L2PHIB11 => return "L1PHIC12_L2PHIB11";
       when L5PHID15_L6PHID27 => return "L5PHID15_L6PHID27";
       when L1PHIF24_L2PHIC23 => return "L1PHIF24_L2PHIC23";
       when L1PHIB8_L2PHIA6 => return "L1PHIB8_L2PHIA6";
       when L1PHIG25_L2PHID27 => return "L1PHIG25_L2PHID27";
       when L2PHII4_L3PHII3 => return "L2PHII4_L3PHII3";
       when L1PHIC9_L2PHIA7 => return "L1PHIC9_L2PHIA7";
       when L3PHID15_L4PHID32 => return "L3PHID15_L4PHID32";
       when L1PHIA4_L2PHIA4 => return "L1PHIA4_L2PHIA4";
       when L1PHIA3_L2PHIA4 => return "L1PHIA3_L2PHIA4";
       when L3PHID16_L4PHID30 => return "L3PHID16_L4PHID30";
       when L1PHIG27_L2PHID29 => return "L1PHIG27_L2PHID29";
       when L5PHID16_L6PHID28 => return "L5PHID16_L6PHID28";
       when L5PHIA4_L6PHIA4 => return "L5PHIA4_L6PHIA4";
       when L3PHIC10_L4PHIC20 => return "L3PHIC10_L4PHIC20";
       when L3PHIC10_L4PHIC18 => return "L3PHIC10_L4PHIC18";
       when L1PHIH32_L2PHID30 => return "L1PHIH32_L2PHID30";
       when L1PHIF22_L2PHIC23 => return "L1PHIF22_L2PHIC23";
       when L5PHIC11_L6PHIC20 => return "L5PHIC11_L6PHIC20";
       when L1PHIC9_L2PHIB11 => return "L1PHIC9_L2PHIB11";
       when L1PHIF23_L2PHIC24 => return "L1PHIF23_L2PHIC24";
       when L5PHID13_L6PHIC23 => return "L5PHID13_L6PHIC23";
       when L1PHID13_L2PHIB13 => return "L1PHID13_L2PHIB13";
       when L5PHID14_L6PHIC24 => return "L5PHID14_L6PHIC24";
       when L1PHIF21_L2PHIC23 => return "L1PHIF21_L2PHIC23";
       when L1PHIG28_L2PHID27 => return "L1PHIG28_L2PHID27";
       when L1PHIE17_L2PHIB15 => return "L1PHIE17_L2PHIB15";
       when L1PHIE18_L2PHIC17 => return "L1PHIE18_L2PHIC17";
       when L5PHIB6_L6PHIB9 => return "L5PHIB6_L6PHIB9";
       when L5PHIB8_L6PHIB16 => return "L5PHIB8_L6PHIB16";
       when L1PHIF23_L2PHIC23 => return "L1PHIF23_L2PHIC23";
       when L1PHIB5_L2PHIA7 => return "L1PHIB5_L2PHIA7";
       when L1PHIH29_L2PHID28 => return "L1PHIH29_L2PHID28";
       when L5PHIC12_L6PHIC22 => return "L5PHIC12_L6PHIC22";
       when L2PHIK11_L3PHIK10 => return "L2PHIK11_L3PHIK10";
       when L5PHID13_L6PHID26 => return "L5PHID13_L6PHID26";
       when L5PHID15_L6PHID28 => return "L5PHID15_L6PHID28";
       when L1PHID14_L2PHIB14 => return "L1PHID14_L2PHIB14";
       when L2PHII2_L3PHII2 => return "L2PHII2_L3PHII2";
       when L2PHIK11_L3PHIK11 => return "L2PHIK11_L3PHIK11";
       when L1PHID15_L2PHIB14 => return "L1PHID15_L2PHIB14";
       when L5PHIC10_L6PHIC23 => return "L5PHIC10_L6PHIC23";
       when L5PHIC11_L6PHID25 => return "L5PHIC11_L6PHID25";
       when L1PHIA1_L2PHIA2 => return "L1PHIA1_L2PHIA2";
       when L5PHID13_L6PHIC24 => return "L5PHID13_L6PHIC24";
       when L1PHID13_L2PHIB12 => return "L1PHID13_L2PHIB12";
       when L3PHIC9_L4PHIC18 => return "L3PHIC9_L4PHIC18";
       when L5PHID15_L6PHID31 => return "L5PHID15_L6PHID31";
       when L1PHIE18_L2PHIC18 => return "L1PHIE18_L2PHIC18";
       when L5PHIB8_L6PHIC17 => return "L5PHIB8_L6PHIC17";
       when L1PHIE18_L2PHIC19 => return "L1PHIE18_L2PHIC19";
       when L1PHIC11_L2PHIB12 => return "L1PHIC11_L2PHIB12";
       when L2PHII3_L3PHII4 => return "L2PHII3_L3PHII4";
       when L5PHIC9_L6PHIC21 => return "L5PHIC9_L6PHIC21";
       when L1PHIG25_L2PHID25 => return "L1PHIG25_L2PHID25";
       when L1PHIB7_L2PHIA7 => return "L1PHIB7_L2PHIA7";
       when L5PHID15_L6PHID30 => return "L5PHID15_L6PHID30";
       when L2PHIJ7_L3PHIJ7 => return "L2PHIJ7_L3PHIJ7";
       when L5PHID13_L6PHID25 => return "L5PHID13_L6PHID25";
       when L2PHIK9_L3PHIK9 => return "L2PHIK9_L3PHIK9";
       when L1PHIC12_L2PHIB13 => return "L1PHIC12_L2PHIB13";
       when L1PHID14_L2PHIB12 => return "L1PHID14_L2PHIB12";
       when L1PHIG25_L2PHIC24 => return "L1PHIG25_L2PHIC24";
       when L5PHIB7_L6PHIB10 => return "L5PHIB7_L6PHIB10";
       when L3PHID14_L4PHID28 => return "L3PHID14_L4PHID28";
       when L1PHIF23_L2PHIC21 => return "L1PHIF23_L2PHIC21";
       when L5PHID13_L6PHIC22 => return "L5PHID13_L6PHIC22";
       when L2PHIK9_L3PHIK10 => return "L2PHIK9_L3PHIK10";
       when L5PHIA4_L6PHIB11 => return "L5PHIA4_L6PHIB11";
       when L1PHIG27_L2PHID27 => return "L1PHIG27_L2PHID27";
       when L1PHID14_L2PHIB13 => return "L1PHID14_L2PHIB13";
       when L5PHIA4_L6PHIB9 => return "L5PHIA4_L6PHIB9";
       when L3PHID13_L4PHIC24 => return "L3PHID13_L4PHIC24";
       when L5PHIB5_L6PHIB9 => return "L5PHIB5_L6PHIB9";
       when L5PHIA1_L6PHIA4 => return "L5PHIA1_L6PHIA4";
       when L1PHIB7_L2PHIA5 => return "L1PHIB7_L2PHIA5";
       when L5PHIA2_L6PHIA2 => return "L5PHIA2_L6PHIA2";
       when L5PHIC9_L6PHIC19 => return "L5PHIC9_L6PHIC19";
       when L1PHIH30_L2PHID31 => return "L1PHIH30_L2PHID31";
       when L1PHIG28_L2PHID28 => return "L1PHIG28_L2PHID28";
       when L5PHID13_L6PHID28 => return "L5PHID13_L6PHID28";
       when L1PHIG26_L2PHID25 => return "L1PHIG26_L2PHID25";
       when L5PHIB5_L6PHIA7 => return "L5PHIB5_L6PHIA7";
       when L1PHIE19_L2PHIC21 => return "L1PHIE19_L2PHIC21";
       when L3PHIB7_L4PHIB14 => return "L3PHIB7_L4PHIB14";
       when L2PHIK10_L3PHIK9 => return "L2PHIK10_L3PHIK9";
       when L3PHID16_L4PHID31 => return "L3PHID16_L4PHID31";
       when L5PHIA3_L6PHIA2 => return "L5PHIA3_L6PHIA2";
       when L3PHIA3_L4PHIA6 => return "L3PHIA3_L4PHIA6";
       when L1PHIH30_L2PHID28 => return "L1PHIH30_L2PHID28";
       when L3PHIB7_L4PHIB12 => return "L3PHIB7_L4PHIB12";
       when L5PHIA1_L6PHIA1 => return "L5PHIA1_L6PHIA1";
       when L5PHIA3_L6PHIA4 => return "L5PHIA3_L6PHIA4";
       when L1PHIC9_L2PHIB10 => return "L1PHIC9_L2PHIB10";
       when L3PHID13_L4PHID28 => return "L3PHID13_L4PHID28";
       when L1PHIH32_L2PHID31 => return "L1PHIH32_L2PHID31";
       when L5PHIB7_L6PHIC17 => return "L5PHIB7_L6PHIC17";
       when L1PHIA3_L2PHIA1 => return "L1PHIA3_L2PHIA1";
       when L2PHII2_L3PHII1 => return "L2PHII2_L3PHII1";
       when L1PHIC12_L2PHIB10 => return "L1PHIC12_L2PHIB10";
       when L2PHIJ7_L3PHIJ6 => return "L2PHIJ7_L3PHIJ6";
       when L1PHIE17_L2PHIC18 => return "L1PHIE17_L2PHIC18";
       when L3PHID15_L4PHID29 => return "L3PHID15_L4PHID29";
       when L2PHIK10_L3PHIK11 => return "L2PHIK10_L3PHIK11";
       when L5PHIA2_L6PHIA7 => return "L5PHIA2_L6PHIA7";
       when L1PHIB5_L2PHIA3 => return "L1PHIB5_L2PHIA3";
       when L1PHIH30_L2PHID32 => return "L1PHIH30_L2PHID32";
       when L3PHIC12_L4PHID26 => return "L3PHIC12_L4PHID26";
       when L3PHIB6_L4PHIB11 => return "L3PHIB6_L4PHIB11";
       when L2PHIL13_L3PHIL14 => return "L2PHIL13_L3PHIL14";
       when L1PHIE19_L2PHIC18 => return "L1PHIE19_L2PHIC18";
       when L1PHIB6_L2PHIA6 => return "L1PHIB6_L2PHIA6";
       when L3PHIC10_L4PHIC19 => return "L3PHIC10_L4PHIC19";
       when L1PHIA2_L2PHIA1 => return "L1PHIA2_L2PHIA1";
       when L1PHIG26_L2PHIC24 => return "L1PHIG26_L2PHIC24";
       when L2PHIJ5_L3PHII4 => return "L2PHIJ5_L3PHII4";
       when L3PHID15_L4PHID31 => return "L3PHID15_L4PHID31";
       when L5PHIB7_L6PHIB11 => return "L5PHIB7_L6PHIB11";
       when L2PHIK11_L3PHIK12 => return "L2PHIK11_L3PHIK12";
       when L3PHIB8_L4PHIB13 => return "L3PHIB8_L4PHIB13";
       when L5PHIB7_L6PHIB13 => return "L5PHIB7_L6PHIB13";
       when L5PHIC10_L6PHIC22 => return "L5PHIC10_L6PHIC22";
       when L3PHIB6_L4PHIB9 => return "L3PHIB6_L4PHIB9";
       when L3PHID16_L4PHID32 => return "L3PHID16_L4PHID32";
       when L5PHIC10_L6PHIB16 => return "L5PHIC10_L6PHIB16";
       when L3PHIA2_L4PHIA3 => return "L3PHIA2_L4PHIA3";
       when L2PHIJ8_L3PHIK9 => return "L2PHIJ8_L3PHIK9";
       when L1PHIC9_L2PHIA8 => return "L1PHIC9_L2PHIA8";
       when L5PHIC10_L6PHIC17 => return "L5PHIC10_L6PHIC17";
       when L3PHIC9_L4PHIC20 => return "L3PHIC9_L4PHIC20";
       when L3PHIB7_L4PHIB13 => return "L3PHIB7_L4PHIB13";
       when L5PHIB7_L6PHIB12 => return "L5PHIB7_L6PHIB12";
       when L5PHIA3_L6PHIB9 => return "L5PHIA3_L6PHIB9";
       when L5PHIA3_L6PHIA7 => return "L5PHIA3_L6PHIA7";
       when L1PHIH31_L2PHID32 => return "L1PHIH31_L2PHID32";
       when L5PHIC9_L6PHIB16 => return "L5PHIC9_L6PHIB16";
       when L1PHIA3_L2PHIA5 => return "L1PHIA3_L2PHIA5";
       when L1PHIF24_L2PHID25 => return "L1PHIF24_L2PHID25";
       when L3PHID16_L4PHID29 => return "L3PHID16_L4PHID29";
       when L3PHIB8_L4PHIC18 => return "L3PHIB8_L4PHIC18";
       when L1PHID15_L2PHIB15 => return "L1PHID15_L2PHIB15";
       when L3PHIB5_L4PHIB11 => return "L3PHIB5_L4PHIB11";
       when L1PHIH31_L2PHID31 => return "L1PHIH31_L2PHID31";
       when L5PHIA4_L6PHIB10 => return "L5PHIA4_L6PHIB10";
       when L3PHIC11_L4PHIC23 => return "L3PHIC11_L4PHIC23";
       when L3PHIA2_L4PHIA6 => return "L3PHIA2_L4PHIA6";
       when L1PHID14_L2PHIB15 => return "L1PHID14_L2PHIB15";
       when L1PHID13_L2PHIB11 => return "L1PHID13_L2PHIB11";
       when L3PHIB7_L4PHIB16 => return "L3PHIB7_L4PHIB16";
       when L1PHIE19_L2PHIC19 => return "L1PHIE19_L2PHIC19";
       when L5PHIB5_L6PHIA6 => return "L5PHIB5_L6PHIA6";
       when L3PHID14_L4PHID26 => return "L3PHID14_L4PHID26";
       when L1PHIB7_L2PHIA8 => return "L1PHIB7_L2PHIA8";
       when L1PHIC10_L2PHIB12 => return "L1PHIC10_L2PHIB12";
       when L3PHIC10_L4PHIC17 => return "L3PHIC10_L4PHIC17";
       when L1PHIG26_L2PHID26 => return "L1PHIG26_L2PHID26";
       when L5PHIC9_L6PHIC20 => return "L5PHIC9_L6PHIC20";
       when L5PHIC9_L6PHIB14 => return "L5PHIC9_L6PHIB14";
       when L5PHID16_L6PHID30 => return "L5PHID16_L6PHID30";
       when L1PHIB8_L2PHIB9 => return "L1PHIB8_L2PHIB9";
       when L1PHIE20_L2PHIC18 => return "L1PHIE20_L2PHIC18";
       when L3PHIA3_L4PHIA8 => return "L3PHIA3_L4PHIA8";
       when L3PHIC11_L4PHIC22 => return "L3PHIC11_L4PHIC22";
       when L1PHIH29_L2PHID31 => return "L1PHIH29_L2PHID31";
       when L3PHIB8_L4PHIC17 => return "L3PHIB8_L4PHIC17";
       when L1PHIA4_L2PHIA2 => return "L1PHIA4_L2PHIA2";
       when L3PHID15_L4PHID28 => return "L3PHID15_L4PHID28";
       when L1PHIF22_L2PHIC20 => return "L1PHIF22_L2PHIC20";
       when L1PHIE17_L2PHIC19 => return "L1PHIE17_L2PHIC19";
       when L5PHIB6_L6PHIB14 => return "L5PHIB6_L6PHIB14";
       when L1PHIF22_L2PHIC22 => return "L1PHIF22_L2PHIC22";
       when L2PHIJ6_L3PHIJ7 => return "L2PHIJ6_L3PHIJ7";
       when L1PHIH30_L2PHID29 => return "L1PHIH30_L2PHID29";
       when L5PHIA2_L6PHIA6 => return "L5PHIA2_L6PHIA6";
       when L5PHIB5_L6PHIB13 => return "L5PHIB5_L6PHIB13";
       when L5PHIA4_L6PHIA7 => return "L5PHIA4_L6PHIA7";
       when L5PHIB5_L6PHIB11 => return "L5PHIB5_L6PHIB11";
       when L2PHIL16_L3PHIL16 => return "L2PHIL16_L3PHIL16";
       when L5PHIC11_L6PHIC21 => return "L5PHIC11_L6PHIC21";
       when L3PHIA4_L4PHIB9 => return "L3PHIA4_L4PHIB9";
       when L5PHID14_L6PHID25 => return "L5PHID14_L6PHID25";
       when L5PHIC10_L6PHIC19 => return "L5PHIC10_L6PHIC19";
       when L5PHID14_L6PHID29 => return "L5PHID14_L6PHID29";
       when L2PHIL16_L3PHIL15 => return "L2PHIL16_L3PHIL15";
       when L1PHIC11_L2PHIB10 => return "L1PHIC11_L2PHIB10";
       when L1PHID15_L2PHIB16 => return "L1PHID15_L2PHIB16";
       when L1PHIG27_L2PHID25 => return "L1PHIG27_L2PHID25";
       when L3PHIB5_L4PHIB9 => return "L3PHIB5_L4PHIB9";
       when L3PHID13_L4PHID27 => return "L3PHID13_L4PHID27";
       when L3PHIB6_L4PHIB14 => return "L3PHIB6_L4PHIB14";
       when L5PHID14_L6PHID27 => return "L5PHID14_L6PHID27";
       when L3PHIC11_L4PHIC19 => return "L3PHIC11_L4PHIC19";
       when L5PHIC12_L6PHID26 => return "L5PHIC12_L6PHID26";
       when L1PHIE20_L2PHIC21 => return "L1PHIE20_L2PHIC21";
       when L1PHIB8_L2PHIA8 => return "L1PHIB8_L2PHIA8";
       when L2PHIJ8_L3PHIJ7 => return "L2PHIJ8_L3PHIJ7";
       when L1PHIF21_L2PHIC19 => return "L1PHIF21_L2PHIC19";
       when L2PHIK9_L3PHIJ8 => return "L2PHIK9_L3PHIJ8";
       when L2PHIL13_L3PHIK12 => return "L2PHIL13_L3PHIK12";
       when L3PHIC9_L4PHIB16 => return "L3PHIC9_L4PHIB16";
       when L5PHIC11_L6PHIC22 => return "L5PHIC11_L6PHIC22";
       when L3PHIA1_L4PHIA2 => return "L3PHIA1_L4PHIA2";
       when L1PHIA3_L2PHIA3 => return "L1PHIA3_L2PHIA3";
       when L2PHIL14_L3PHIL13 => return "L2PHIL14_L3PHIL13";
       when L3PHIB5_L4PHIB10 => return "L3PHIB5_L4PHIB10";
       when L3PHID15_L4PHID30 => return "L3PHID15_L4PHID30";
       when L1PHIB5_L2PHIA5 => return "L1PHIB5_L2PHIA5";
       when L1PHID16_L2PHIC18 => return "L1PHID16_L2PHIC18";
       when L1PHIH31_L2PHID30 => return "L1PHIH31_L2PHID30";
       when L1PHIA2_L2PHIA4 => return "L1PHIA2_L2PHIA4";
       when L5PHID15_L6PHID32 => return "L5PHID15_L6PHID32";
       when L3PHID14_L4PHID27 => return "L3PHID14_L4PHID27";
       when L2PHIJ7_L3PHIJ8 => return "L2PHIJ7_L3PHIJ8";
       when L5PHIA1_L6PHIA3 => return "L5PHIA1_L6PHIA3";
       when L1PHIC10_L2PHIA8 => return "L1PHIC10_L2PHIA8";
       when L1PHIB6_L2PHIA7 => return "L1PHIB6_L2PHIA7";
       when L5PHIA2_L6PHIA1 => return "L5PHIA2_L6PHIA1";
       when L5PHIA4_L6PHIA5 => return "L5PHIA4_L6PHIA5";
       when L1PHIF24_L2PHID26 => return "L1PHIF24_L2PHID26";
       when L2PHII1_L3PHII1 => return "L2PHII1_L3PHII1";
       when L5PHIA2_L6PHIA3 => return "L5PHIA2_L6PHIA3";
       when L5PHIB5_L6PHIB10 => return "L5PHIB5_L6PHIB10";
       when L3PHIA4_L4PHIB10 => return "L3PHIA4_L4PHIB10";
       when L3PHIC10_L4PHIC22 => return "L3PHIC10_L4PHIC22";
       when L3PHIA2_L4PHIA4 => return "L3PHIA2_L4PHIA4";
       when L2PHIL15_L3PHIL15 => return "L2PHIL15_L3PHIL15";
       when L1PHIF21_L2PHIC20 => return "L1PHIF21_L2PHIC20";
       when L1PHIA1_L2PHIA1 => return "L1PHIA1_L2PHIA1";
       when L3PHIB7_L4PHIB15 => return "L3PHIB7_L4PHIB15";
       when L1PHIE17_L2PHIC17 => return "L1PHIE17_L2PHIC17";
       when L5PHIB6_L6PHIA8 => return "L5PHIB6_L6PHIA8";
       when L1PHIF22_L2PHIC21 => return "L1PHIF22_L2PHIC21";
       when L1PHIE20_L2PHIC22 => return "L1PHIE20_L2PHIC22";
       when L5PHIC9_L6PHIB15 => return "L5PHIC9_L6PHIB15";
       when L1PHIG27_L2PHID26 => return "L1PHIG27_L2PHID26";
       when L5PHIC10_L6PHIC21 => return "L5PHIC10_L6PHIC21";
       when L1PHIG28_L2PHID26 => return "L1PHIG28_L2PHID26";
       when L2PHIJ8_L3PHIJ8 => return "L2PHIJ8_L3PHIJ8";
       when L5PHIC11_L6PHIC19 => return "L5PHIC11_L6PHIC19";
       when L1PHIC10_L2PHIB10 => return "L1PHIC10_L2PHIB10";
       when L2PHIJ6_L3PHIJ5 => return "L2PHIJ6_L3PHIJ5";
       when L1PHIG25_L2PHIC23 => return "L1PHIG25_L2PHIC23";
       when L1PHID16_L2PHIB16 => return "L1PHID16_L2PHIB16";
       when L3PHIB6_L4PHIB12 => return "L3PHIB6_L4PHIB12";
       when L3PHIB8_L4PHIB15 => return "L3PHIB8_L4PHIB15";
       when L1PHIC11_L2PHIB9 => return "L1PHIC11_L2PHIB9";
       when L3PHIC9_L4PHIB15 => return "L3PHIC9_L4PHIB15";
       when L1PHIE20_L2PHIC20 => return "L1PHIE20_L2PHIC20";
       when L1PHIB6_L2PHIA5 => return "L1PHIB6_L2PHIA5";
       when L1PHIC11_L2PHIB13 => return "L1PHIC11_L2PHIB13";
       when L1PHIC11_L2PHIB11 => return "L1PHIC11_L2PHIB11";
       when L5PHIB5_L6PHIA8 => return "L5PHIB5_L6PHIA8";
       when L2PHIL15_L3PHIL16 => return "L2PHIL15_L3PHIL16";
       when L3PHID14_L4PHID30 => return "L3PHID14_L4PHID30";
       when L1PHIB6_L2PHIA8 => return "L1PHIB6_L2PHIA8";
       when L1PHID16_L2PHIC17 => return "L1PHID16_L2PHIC17";
       when L1PHID15_L2PHIB13 => return "L1PHID15_L2PHIB13";
       when L1PHIF22_L2PHIC24 => return "L1PHIF22_L2PHIC24";
       when L1PHIB7_L2PHIA6 => return "L1PHIB7_L2PHIA6";
       when L3PHID15_L4PHID27 => return "L3PHID15_L4PHID27";
       when L1PHIH29_L2PHID27 => return "L1PHIH29_L2PHID27";
       when L5PHIB8_L6PHIB15 => return "L5PHIB8_L6PHIB15";
       when L3PHIB5_L4PHIB12 => return "L3PHIB5_L4PHIB12";
       when L2PHIJ6_L3PHIJ6 => return "L2PHIJ6_L3PHIJ6";
       when L5PHIA1_L6PHIA5 => return "L5PHIA1_L6PHIA5";
       when L1PHIE20_L2PHIC19 => return "L1PHIE20_L2PHIC19";
       when L3PHIC12_L4PHID25 => return "L3PHIC12_L4PHID25";
       when L5PHIB6_L6PHIB15 => return "L5PHIB6_L6PHIB15";
       when L1PHID13_L2PHIB14 => return "L1PHID13_L2PHIB14";
       when L5PHIB7_L6PHIB15 => return "L5PHIB7_L6PHIB15";
       when L2PHIL14_L3PHIL14 => return "L2PHIL14_L3PHIL14";
       when L5PHIC11_L6PHIC24 => return "L5PHIC11_L6PHIC24";
       when L2PHII2_L3PHII3 => return "L2PHII2_L3PHII3";
       when L1PHIB8_L2PHIA7 => return "L1PHIB8_L2PHIA7";
       when L1PHID13_L2PHIB15 => return "L1PHID13_L2PHIB15";
       when L5PHIC9_L6PHIC17 => return "L5PHIC9_L6PHIC17";
       when L5PHID15_L6PHID26 => return "L5PHID15_L6PHID26";
       when L5PHIA2_L6PHIA4 => return "L5PHIA2_L6PHIA4";
       when L3PHIB8_L4PHIB16 => return "L3PHIB8_L4PHIB16";
       when L2PHIL13_L3PHIL13 => return "L2PHIL13_L3PHIL13";
       when L1PHIA2_L2PHIA3 => return "L1PHIA2_L2PHIA3";
       when L3PHIC12_L4PHIC24 => return "L3PHIC12_L4PHIC24";
       when L5PHIB6_L6PHIB11 => return "L5PHIB6_L6PHIB11";
       when L1PHIB5_L2PHIA4 => return "L1PHIB5_L2PHIA4";
       when L5PHIA3_L6PHIA8 => return "L5PHIA3_L6PHIA8";
       when L5PHIB7_L6PHIB14 => return "L5PHIB7_L6PHIB14";
       when L2PHIK12_L3PHIK11 => return "L2PHIK12_L3PHIK11";
       when L1PHIH29_L2PHID30 => return "L1PHIH29_L2PHID30";
       when L3PHID13_L4PHIC23 => return "L3PHID13_L4PHIC23";
       when L1PHIC12_L2PHIB14 => return "L1PHIC12_L2PHIB14";
       when L5PHID14_L6PHID30 => return "L5PHID14_L6PHID30";
       when L1PHIH29_L2PHID29 => return "L1PHIH29_L2PHID29";
       when L1PHIF23_L2PHIC22 => return "L1PHIF23_L2PHIC22";
       when L5PHID16_L6PHID31 => return "L5PHID16_L6PHID31";
       when L2PHII4_L3PHIJ5 => return "L2PHII4_L3PHIJ5";
       when L5PHIA3_L6PHIA3 => return "L5PHIA3_L6PHIA3";
       when L3PHIB6_L4PHIB13 => return "L3PHIB6_L4PHIB13";
       when L1PHID14_L2PHIB16 => return "L1PHID14_L2PHIB16";
       when L5PHIC9_L6PHIC18 => return "L5PHIC9_L6PHIC18";
       when L1PHIB6_L2PHIA4 => return "L1PHIB6_L2PHIA4";
       when L5PHIC12_L6PHID25 => return "L5PHIC12_L6PHID25";
       when L5PHIB7_L6PHIB16 => return "L5PHIB7_L6PHIB16";
       when L1PHIA4_L2PHIA3 => return "L1PHIA4_L2PHIA3";
       when L3PHIA2_L4PHIA5 => return "L3PHIA2_L4PHIA5";
       when L5PHIA2_L6PHIA5 => return "L5PHIA2_L6PHIA5";
       when L2PHIJ5_L3PHIJ6 => return "L2PHIJ5_L3PHIJ6";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_TPROJ_60) return string is
  begin
    case val is
       when L5L6C_L1PHIC => return "L5L6C_L1PHIC";
       when L2L3C_L1PHIE => return "L2L3C_L1PHIE";
       when L5L6A_L2PHIA => return "L5L6A_L2PHIA";
       when L5L6A_L1PHIA => return "L5L6A_L1PHIA";
       when L3L4C_L2PHIC => return "L3L4C_L2PHIC";
       when L5L6B_L2PHIB => return "L5L6B_L2PHIB";
       when L3L4B_L1PHIE => return "L3L4B_L1PHIE";
       when L3L4D_L2PHID => return "L3L4D_L2PHID";
       when L3L4C_L1PHIG => return "L3L4C_L1PHIG";
       when L1L2K_L3PHID => return "L1L2K_L3PHID";
       when L3L4B_L1PHID => return "L3L4B_L1PHID";
       when L5L6C_L1PHIF => return "L5L6C_L1PHIF";
       when L5L6C_L1PHIE => return "L5L6C_L1PHIE";
       when L3L4B_L2PHIA => return "L3L4B_L2PHIA";
       when L2L3C_L1PHIF => return "L2L3C_L1PHIF";
       when L1L2J_L3PHID => return "L1L2J_L3PHID";
       when L5L6B_L1PHID => return "L5L6B_L1PHID";
       when L1L2J_L3PHIC => return "L1L2J_L3PHIC";
       when L1L2I_L3PHID => return "L1L2I_L3PHID";
       when L1L2E_L3PHIB => return "L1L2E_L3PHIB";
       when L2L3A_L1PHIC => return "L2L3A_L1PHIC";
       when L5L6B_L1PHIF => return "L5L6B_L1PHIF";
       when L5L6A_L1PHID => return "L5L6A_L1PHID";
       when L3L4C_L1PHIE => return "L3L4C_L1PHIE";
       when L5L6C_L2PHID => return "L5L6C_L2PHID";
       when L1L2G_L3PHIC => return "L1L2G_L3PHIC";
       when L3L4B_L2PHIC => return "L3L4B_L2PHIC";
       when L3L4B_L1PHIC => return "L3L4B_L1PHIC";
       when L2L3D_L1PHIH => return "L2L3D_L1PHIH";
       when L5L6B_L1PHIC => return "L5L6B_L1PHIC";
       when L1L2F_L3PHIB => return "L1L2F_L3PHIB";
       when L1L2D_L3PHIA => return "L1L2D_L3PHIA";
       when L3L4D_L2PHIC => return "L3L4D_L2PHIC";
       when L3L4A_L1PHIB => return "L3L4A_L1PHIB";
       when L1L2F_L3PHIC => return "L1L2F_L3PHIC";
       when L1L2I_L3PHIC => return "L1L2I_L3PHIC";
       when L2L3D_L1PHIG => return "L2L3D_L1PHIG";
       when L3L4A_L1PHIC => return "L3L4A_L1PHIC";
       when L3L4A_L2PHIB => return "L3L4A_L2PHIB";
       when L1L2H_L3PHIC => return "L1L2H_L3PHIC";
       when L5L6A_L1PHIC => return "L5L6A_L1PHIC";
       when L5L6A_L3PHIA => return "L5L6A_L3PHIA";
       when L5L6D_L2PHID => return "L5L6D_L2PHID";
       when L5L6D_L1PHIE => return "L5L6D_L1PHIE";
       when L5L6D_L1PHIH => return "L5L6D_L1PHIH";
       when L5L6B_L1PHIB => return "L5L6B_L1PHIB";
       when L1L2C_L3PHIA => return "L1L2C_L3PHIA";
       when L5L6B_L2PHIC => return "L5L6B_L2PHIC";
       when L3L4B_L1PHIB => return "L3L4B_L1PHIB";
       when L2L3A_L1PHIB => return "L2L3A_L1PHIB";
       when L2L3B_L1PHIC => return "L2L3B_L1PHIC";
       when L5L6B_L3PHIA => return "L5L6B_L3PHIA";
       when L2L3B_L1PHIE => return "L2L3B_L1PHIE";
       when L3L4D_L1PHIH => return "L3L4D_L1PHIH";
       when L1L2A_L3PHIA => return "L1L2A_L3PHIA";
       when L2L3C_L1PHID => return "L2L3C_L1PHID";
       when L3L4A_L1PHIA => return "L3L4A_L1PHIA";
       when L5L6D_L1PHIF => return "L5L6D_L1PHIF";
       when L2L3C_L1PHIG => return "L2L3C_L1PHIG";
       when L1L2B_L3PHIB => return "L1L2B_L3PHIB";
       when L5L6B_L3PHIC => return "L5L6B_L3PHIC";
       when L2L3A_L1PHIA => return "L2L3A_L1PHIA";
       when L5L6D_L3PHIC => return "L5L6D_L3PHIC";
       when L5L6B_L2PHIA => return "L5L6B_L2PHIA";
       when L1L2G_L3PHIB => return "L1L2G_L3PHIB";
       when L3L4B_L2PHIB => return "L3L4B_L2PHIB";
       when L1L2L_L3PHID => return "L1L2L_L3PHID";
       when L5L6B_L3PHIB => return "L5L6B_L3PHIB";
       when L5L6A_L3PHIB => return "L5L6A_L3PHIB";
       when L5L6A_L1PHIB => return "L5L6A_L1PHIB";
       when L5L6C_L3PHIB => return "L5L6C_L3PHIB";
       when L5L6D_L3PHID => return "L5L6D_L3PHID";
       when L2L3D_L1PHIF => return "L2L3D_L1PHIF";
       when L5L6C_L3PHID => return "L5L6C_L3PHID";
       when L5L6B_L1PHIE => return "L5L6B_L1PHIE";
       when L5L6C_L3PHIC => return "L5L6C_L3PHIC";
       when L1L2B_L3PHIA => return "L1L2B_L3PHIA";
       when L5L6C_L1PHID => return "L5L6C_L1PHID";
       when L3L4C_L1PHIF => return "L3L4C_L1PHIF";
       when L1L2D_L3PHIB => return "L1L2D_L3PHIB";
       when L1L2C_L3PHIB => return "L1L2C_L3PHIB";
       when L3L4C_L2PHIB => return "L3L4C_L2PHIB";
       when L5L6C_L2PHIC => return "L5L6C_L2PHIC";
       when L3L4C_L2PHID => return "L3L4C_L2PHID";
       when L2L3B_L1PHID => return "L2L3B_L1PHID";
       when L5L6C_L2PHIB => return "L5L6C_L2PHIB";
       when L3L4A_L2PHIA => return "L3L4A_L2PHIA";
       when L3L4D_L1PHIG => return "L3L4D_L1PHIG";
       when L5L6D_L2PHIC => return "L5L6D_L2PHIC";
       when L5L6C_L1PHIG => return "L5L6C_L1PHIG";
       when L5L6D_L1PHIG => return "L5L6D_L1PHIG";
       when L3L4C_L1PHID => return "L3L4C_L1PHID";
       when L5L6A_L2PHIB => return "L5L6A_L2PHIB";
       when L3L4D_L1PHIF => return "L3L4D_L1PHIF";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_TPROJ_58) return string is
  begin
    case val is
       when L2L3C_L5PHIB => return "L2L3C_L5PHIB";
       when L1L2E_L5PHIC => return "L1L2E_L5PHIC";
       when L1L2H_L6PHIC => return "L1L2H_L6PHIC";
       when L3L4B_L5PHIA => return "L3L4B_L5PHIA";
       when L3L4C_L5PHIB => return "L3L4C_L5PHIB";
       when L1L2L_L6PHIC => return "L1L2L_L6PHIC";
       when L1L2H_L4PHIB => return "L1L2H_L4PHIB";
       when L1L2H_L5PHID => return "L1L2H_L5PHID";
       when L1L2L_L4PHID => return "L1L2L_L4PHID";
       when L2L3C_L5PHID => return "L2L3C_L5PHID";
       when L1L2H_L6PHID => return "L1L2H_L6PHID";
       when L1L2E_L6PHIB => return "L1L2E_L6PHIB";
       when L1L2J_L6PHID => return "L1L2J_L6PHID";
       when L1L2L_L5PHID => return "L1L2L_L5PHID";
       when L1L2K_L4PHID => return "L1L2K_L4PHID";
       when L1L2H_L4PHIC => return "L1L2H_L4PHIC";
       when L3L4B_L5PHIC => return "L3L4B_L5PHIC";
       when L1L2K_L4PHIC => return "L1L2K_L4PHIC";
       when L1L2G_L4PHIC => return "L1L2G_L4PHIC";
       when L3L4D_L6PHIC => return "L3L4D_L6PHIC";
       when L5L6A_L4PHIA => return "L5L6A_L4PHIA";
       when L3L4C_L5PHID => return "L3L4C_L5PHID";
       when L1L2A_L5PHIB => return "L1L2A_L5PHIB";
       when L2L3B_L5PHIB => return "L2L3B_L5PHIB";
       when L1L2C_L6PHIB => return "L1L2C_L6PHIB";
       when L3L4D_L6PHID => return "L3L4D_L6PHID";
       when L5L6A_L4PHIB => return "L5L6A_L4PHIB";
       when L5L6D_L4PHID => return "L5L6D_L4PHID";
       when L1L2G_L6PHID => return "L1L2G_L6PHID";
       when L2L3D_L4PHID => return "L2L3D_L4PHID";
       when L1L2D_L5PHIC => return "L1L2D_L5PHIC";
       when L1L2I_L5PHID => return "L1L2I_L5PHID";
       when L1L2E_L4PHIC => return "L1L2E_L4PHIC";
       when L1L2E_L4PHIA => return "L1L2E_L4PHIA";
       when L2L3B_L4PHIA => return "L2L3B_L4PHIA";
       when L1L2I_L4PHIC => return "L1L2I_L4PHIC";
       when L1L2I_L4PHID => return "L1L2I_L4PHID";
       when L1L2G_L6PHIB => return "L1L2G_L6PHIB";
       when L2L3D_L5PHIC => return "L2L3D_L5PHIC";
       when L1L2F_L5PHIC => return "L1L2F_L5PHIC";
       when L2L3A_L4PHIA => return "L2L3A_L4PHIA";
       when L5L6C_L4PHIB => return "L5L6C_L4PHIB";
       when L1L2B_L5PHIA => return "L1L2B_L5PHIA";
       when L1L2G_L4PHIB => return "L1L2G_L4PHIB";
       when L1L2F_L6PHIA => return "L1L2F_L6PHIA";
       when L1L2H_L5PHIB => return "L1L2H_L5PHIB";
       when L2L3B_L5PHIC => return "L2L3B_L5PHIC";
       when L1L2H_L5PHIC => return "L1L2H_L5PHIC";
       when L1L2J_L5PHID => return "L1L2J_L5PHID";
       when L1L2D_L4PHIA => return "L1L2D_L4PHIA";
       when L1L2D_L6PHIB => return "L1L2D_L6PHIB";
       when L1L2I_L5PHIB => return "L1L2I_L5PHIB";
       when L1L2A_L4PHIA => return "L1L2A_L4PHIA";
       when L1L2D_L6PHIA => return "L1L2D_L6PHIA";
       when L1L2C_L4PHIA => return "L1L2C_L4PHIA";
       when L3L4A_L6PHIA => return "L3L4A_L6PHIA";
       when L1L2A_L6PHIB => return "L1L2A_L6PHIB";
       when L2L3A_L5PHIA => return "L2L3A_L5PHIA";
       when L3L4D_L5PHID => return "L3L4D_L5PHID";
       when L1L2E_L4PHIB => return "L1L2E_L4PHIB";
       when L5L6B_L4PHIC => return "L5L6B_L4PHIC";
       when L2L3D_L5PHID => return "L2L3D_L5PHID";
       when L1L2C_L5PHIA => return "L1L2C_L5PHIA";
       when L1L2I_L6PHID => return "L1L2I_L6PHID";
       when L3L4C_L6PHIB => return "L3L4C_L6PHIB";
       when L3L4C_L6PHIC => return "L3L4C_L6PHIC";
       when L2L3A_L5PHIB => return "L2L3A_L5PHIB";
       when L1L2J_L5PHIC => return "L1L2J_L5PHIC";
       when L1L2B_L4PHIA => return "L1L2B_L4PHIA";
       when L3L4A_L5PHIA => return "L3L4A_L5PHIA";
       when L1L2A_L5PHIA => return "L1L2A_L5PHIA";
       when L3L4B_L6PHIA => return "L3L4B_L6PHIA";
       when L1L2C_L4PHIB => return "L1L2C_L4PHIB";
       when L1L2B_L6PHIB => return "L1L2B_L6PHIB";
       when L1L2B_L4PHIB => return "L1L2B_L4PHIB";
       when L2L3D_L4PHIC => return "L2L3D_L4PHIC";
       when L1L2G_L5PHIC => return "L1L2G_L5PHIC";
       when L1L2E_L6PHIA => return "L1L2E_L6PHIA";
       when L5L6B_L4PHIB => return "L5L6B_L4PHIB";
       when L1L2G_L6PHIC => return "L1L2G_L6PHIC";
       when L3L4B_L5PHIB => return "L3L4B_L5PHIB";
       when L2L3A_L4PHIB => return "L2L3A_L4PHIB";
       when L1L2I_L6PHIC => return "L1L2I_L6PHIC";
       when L1L2C_L6PHIA => return "L1L2C_L6PHIA";
       when L2L3B_L4PHIB => return "L2L3B_L4PHIB";
       when L1L2J_L4PHID => return "L1L2J_L4PHID";
       when L1L2F_L5PHIB => return "L1L2F_L5PHIB";
       when L1L2D_L6PHIC => return "L1L2D_L6PHIC";
       when L1L2K_L6PHIC => return "L1L2K_L6PHIC";
       when L1L2H_L6PHIB => return "L1L2H_L6PHIB";
       when L1L2K_L5PHIC => return "L1L2K_L5PHIC";
       when L3L4C_L6PHID => return "L3L4C_L6PHID";
       when L1L2K_L6PHID => return "L1L2K_L6PHID";
       when L2L3C_L4PHIB => return "L2L3C_L4PHIB";
       when L1L2L_L5PHIC => return "L1L2L_L5PHIC";
       when L5L6C_L4PHIC => return "L5L6C_L4PHIC";
       when L3L4A_L6PHIB => return "L3L4A_L6PHIB";
       when L1L2D_L5PHIA => return "L1L2D_L5PHIA";
       when L1L2F_L4PHIC => return "L1L2F_L4PHIC";
       when L1L2J_L4PHIC => return "L1L2J_L4PHIC";
       when L1L2J_L6PHIC => return "L1L2J_L6PHIC";
       when L1L2E_L5PHIA => return "L1L2E_L5PHIA";
       when L1L2B_L5PHIB => return "L1L2B_L5PHIB";
       when L1L2I_L6PHIB => return "L1L2I_L6PHIB";
       when L2L3C_L4PHIC => return "L2L3C_L4PHIC";
       when L1L2E_L5PHIB => return "L1L2E_L5PHIB";
       when L1L2G_L5PHIB => return "L1L2G_L5PHIB";
       when L3L4C_L5PHIC => return "L3L4C_L5PHIC";
       when L3L4A_L5PHIB => return "L3L4A_L5PHIB";
       when L1L2E_L6PHIC => return "L1L2E_L6PHIC";
       when L1L2C_L5PHIB => return "L1L2C_L5PHIB";
       when L5L6B_L4PHIA => return "L5L6B_L4PHIA";
       when L2L3B_L5PHIA => return "L2L3B_L5PHIA";
       when L2L3C_L4PHID => return "L2L3C_L4PHID";
       when L1L2B_L6PHIA => return "L1L2B_L6PHIA";
       when L1L2I_L5PHIC => return "L1L2I_L5PHIC";
       when L5L6D_L4PHIC => return "L5L6D_L4PHIC";
       when L2L3C_L5PHIC => return "L2L3C_L5PHIC";
       when L1L2H_L4PHID => return "L1L2H_L4PHID";
       when L1L2F_L6PHIC => return "L1L2F_L6PHIC";
       when L1L2F_L6PHIB => return "L1L2F_L6PHIB";
       when L3L4B_L6PHIC => return "L3L4B_L6PHIC";
       when L5L6C_L4PHID => return "L5L6C_L4PHID";
       when L1L2D_L5PHIB => return "L1L2D_L5PHIB";
       when L1L2F_L4PHIB => return "L1L2F_L4PHIB";
       when L1L2K_L5PHID => return "L1L2K_L5PHID";
       when L1L2D_L4PHIB => return "L1L2D_L4PHIB";
       when L2L3B_L4PHIC => return "L2L3B_L4PHIC";
       when L3L4B_L6PHIB => return "L3L4B_L6PHIB";
       when L3L4D_L5PHIC => return "L3L4D_L5PHIC";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_TPAR_70) return string is
  begin
    case val is
       when L1L2F => return "L1L2F";
       when L1L2I => return "L1L2I";
       when L1L2D => return "L1L2D";
       when L2L3B => return "L2L3B";
       when L3L4D => return "L3L4D";
       when L3L4A => return "L3L4A";
       when L3L4C => return "L3L4C";
       when L5L6C => return "L5L6C";
       when L1L2E => return "L1L2E";
       when L5L6A => return "L5L6A";
       when L2L3D => return "L2L3D";
       when L1L2C => return "L1L2C";
       when L1L2J => return "L1L2J";
       when L5L6B => return "L5L6B";
       when L1L2B => return "L1L2B";
       when L2L3A => return "L2L3A";
       when L1L2K => return "L1L2K";
       when L1L2L => return "L1L2L";
       when L1L2H => return "L1L2H";
       when L2L3C => return "L2L3C";
       when L1L2G => return "L1L2G";
       when L3L4B => return "L3L4B";
       when L5L6D => return "L5L6D";
       when L1L2A => return "L1L2A";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_VMPROJ_24) return string is
  begin
    case val is
       when L4PHIB16 => return "L4PHIB16";
       when L2PHID26 => return "L2PHID26";
       when L4PHID32 => return "L4PHID32";
       when L4PHID25 => return "L4PHID25";
       when L5PHIC22 => return "L5PHIC22";
       when L3PHIC24 => return "L3PHIC24";
       when L4PHIA5 => return "L4PHIA5";
       when L6PHID28 => return "L6PHID28";
       when L6PHIB11 => return "L6PHIB11";
       when L2PHIB10 => return "L2PHIB10";
       when L1PHIA4 => return "L1PHIA4";
       when L3PHIC17 => return "L3PHIC17";
       when L2PHID25 => return "L2PHID25";
       when L6PHID26 => return "L6PHID26";
       when L1PHIC10 => return "L1PHIC10";
       when L2PHID28 => return "L2PHID28";
       when L6PHID31 => return "L6PHID31";
       when L6PHIA3 => return "L6PHIA3";
       when L2PHIC19 => return "L2PHIC19";
       when L1PHID16 => return "L1PHID16";
       when L3PHID26 => return "L3PHID26";
       when L3PHID28 => return "L3PHID28";
       when L4PHIA7 => return "L4PHIA7";
       when L4PHIC19 => return "L4PHIC19";
       when L1PHID14 => return "L1PHID14";
       when L3PHIC21 => return "L3PHIC21";
       when L6PHIA2 => return "L6PHIA2";
       when L5PHIA7 => return "L5PHIA7";
       when L6PHIB13 => return "L6PHIB13";
       when L4PHIA3 => return "L4PHIA3";
       when L4PHIA4 => return "L4PHIA4";
       when L4PHIC24 => return "L4PHIC24";
       when L5PHIB9 => return "L5PHIB9";
       when L3PHIA5 => return "L3PHIA5";
       when L4PHIB12 => return "L4PHIB12";
       when L3PHIC18 => return "L3PHIC18";
       when L5PHIA5 => return "L5PHIA5";
       when L1PHIE19 => return "L1PHIE19";
       when L3PHIC19 => return "L3PHIC19";
       when L3PHIA8 => return "L3PHIA8";
       when L2PHIA7 => return "L2PHIA7";
       when L6PHIB15 => return "L6PHIB15";
       when L5PHIB12 => return "L5PHIB12";
       when L4PHIC20 => return "L4PHIC20";
       when L2PHIB14 => return "L2PHIB14";
       when L1PHIG28 => return "L1PHIG28";
       when L1PHIB5 => return "L1PHIB5";
       when L3PHIB11 => return "L3PHIB11";
       when L6PHIC23 => return "L6PHIC23";
       when L5PHID32 => return "L5PHID32";
       when L2PHIA5 => return "L2PHIA5";
       when L3PHIB16 => return "L3PHIB16";
       when L2PHIB15 => return "L2PHIB15";
       when L5PHIA8 => return "L5PHIA8";
       when L2PHIA3 => return "L2PHIA3";
       when L1PHIH31 => return "L1PHIH31";
       when L1PHIC11 => return "L1PHIC11";
       when L1PHIB6 => return "L1PHIB6";
       when L2PHIB9 => return "L2PHIB9";
       when L1PHIH32 => return "L1PHIH32";
       when L1PHIG27 => return "L1PHIG27";
       when L4PHIB9 => return "L4PHIB9";
       when L2PHIA8 => return "L2PHIA8";
       when L5PHID27 => return "L5PHID27";
       when L6PHIA8 => return "L6PHIA8";
       when L3PHID25 => return "L3PHID25";
       when L5PHIB15 => return "L5PHIB15";
       when L1PHIH29 => return "L1PHIH29";
       when L4PHID30 => return "L4PHID30";
       when L3PHIC22 => return "L3PHIC22";
       when L6PHID29 => return "L6PHID29";
       when L5PHIA4 => return "L5PHIA4";
       when L1PHID15 => return "L1PHID15";
       when L5PHID30 => return "L5PHID30";
       when L4PHID31 => return "L4PHID31";
       when L6PHIC20 => return "L6PHIC20";
       when L6PHIA4 => return "L6PHIA4";
       when L4PHID26 => return "L4PHID26";
       when L5PHIC21 => return "L5PHIC21";
       when L2PHIC23 => return "L2PHIC23";
       when L4PHIA8 => return "L4PHIA8";
       when L5PHID29 => return "L5PHID29";
       when L3PHID29 => return "L3PHID29";
       when L4PHIB14 => return "L4PHIB14";
       when L4PHIA6 => return "L4PHIA6";
       when L3PHIB10 => return "L3PHIB10";
       when L2PHIA1 => return "L2PHIA1";
       when L4PHIB11 => return "L4PHIB11";
       when L5PHIA2 => return "L5PHIA2";
       when L6PHIC17 => return "L6PHIC17";
       when L1PHIA2 => return "L1PHIA2";
       when L3PHID27 => return "L3PHID27";
       when L1PHIF21 => return "L1PHIF21";
       when L6PHIB9 => return "L6PHIB9";
       when L5PHIC17 => return "L5PHIC17";
       when L5PHIA6 => return "L5PHIA6";
       when L1PHIF23 => return "L1PHIF23";
       when L5PHID28 => return "L5PHID28";
       when L1PHIB8 => return "L1PHIB8";
       when L3PHIA1 => return "L3PHIA1";
       when L5PHID26 => return "L5PHID26";
       when L5PHIC20 => return "L5PHIC20";
       when L1PHID13 => return "L1PHID13";
       when L2PHIC18 => return "L2PHIC18";
       when L3PHIA7 => return "L3PHIA7";
       when L6PHIC18 => return "L6PHIC18";
       when L6PHIC21 => return "L6PHIC21";
       when L4PHIC22 => return "L4PHIC22";
       when L2PHID32 => return "L2PHID32";
       when L3PHID32 => return "L3PHID32";
       when L6PHID27 => return "L6PHID27";
       when L1PHIC9 => return "L1PHIC9";
       when L5PHIA3 => return "L5PHIA3";
       when L2PHIB13 => return "L2PHIB13";
       when L2PHIC17 => return "L2PHIC17";
       when L4PHIB15 => return "L4PHIB15";
       when L1PHIA1 => return "L1PHIA1";
       when L6PHIA5 => return "L6PHIA5";
       when L5PHIB10 => return "L5PHIB10";
       when L1PHIC12 => return "L1PHIC12";
       when L4PHIA1 => return "L4PHIA1";
       when L1PHIE17 => return "L1PHIE17";
       when L3PHID31 => return "L3PHID31";
       when L2PHIA6 => return "L2PHIA6";
       when L3PHIA4 => return "L3PHIA4";
       when L2PHIC20 => return "L2PHIC20";
       when L6PHIB16 => return "L6PHIB16";
       when L1PHIB7 => return "L1PHIB7";
       when L2PHID29 => return "L2PHID29";
       when L6PHID32 => return "L6PHID32";
       when L4PHIC21 => return "L4PHIC21";
       when L4PHIB10 => return "L4PHIB10";
       when L3PHIA6 => return "L3PHIA6";
       when L6PHID30 => return "L6PHID30";
       when L3PHIB12 => return "L3PHIB12";
       when L5PHIB14 => return "L5PHIB14";
       when L5PHIC23 => return "L5PHIC23";
       when L5PHIC24 => return "L5PHIC24";
       when L6PHIB10 => return "L6PHIB10";
       when L2PHIC24 => return "L2PHIC24";
       when L4PHID28 => return "L4PHID28";
       when L5PHIA1 => return "L5PHIA1";
       when L6PHIC22 => return "L6PHIC22";
       when L4PHIC17 => return "L4PHIC17";
       when L3PHIB14 => return "L3PHIB14";
       when L5PHID25 => return "L5PHID25";
       when L2PHIA4 => return "L2PHIA4";
       when L5PHIC19 => return "L5PHIC19";
       when L6PHIC24 => return "L6PHIC24";
       when L6PHIB12 => return "L6PHIB12";
       when L4PHIB13 => return "L4PHIB13";
       when L6PHIA1 => return "L6PHIA1";
       when L6PHIA6 => return "L6PHIA6";
       when L2PHID31 => return "L2PHID31";
       when L3PHIB15 => return "L3PHIB15";
       when L4PHID27 => return "L4PHID27";
       when L1PHIA3 => return "L1PHIA3";
       when L2PHIC22 => return "L2PHIC22";
       when L6PHIC19 => return "L6PHIC19";
       when L2PHIA2 => return "L2PHIA2";
       when L1PHIG25 => return "L1PHIG25";
       when L4PHIC23 => return "L4PHIC23";
       when L2PHIC21 => return "L2PHIC21";
       when L6PHIB14 => return "L6PHIB14";
       when L6PHID25 => return "L6PHID25";
       when L1PHIF22 => return "L1PHIF22";
       when L2PHID27 => return "L2PHID27";
       when L4PHIC18 => return "L4PHIC18";
       when L1PHIF24 => return "L1PHIF24";
       when L3PHIB13 => return "L3PHIB13";
       when L1PHIH30 => return "L1PHIH30";
       when L3PHIC20 => return "L3PHIC20";
       when L2PHIB16 => return "L2PHIB16";
       when L2PHIB12 => return "L2PHIB12";
       when L3PHID30 => return "L3PHID30";
       when L1PHIE18 => return "L1PHIE18";
       when L5PHIC18 => return "L5PHIC18";
       when L2PHID30 => return "L2PHID30";
       when L6PHIA7 => return "L6PHIA7";
       when L5PHIB11 => return "L5PHIB11";
       when L3PHIA3 => return "L3PHIA3";
       when L1PHIE20 => return "L1PHIE20";
       when L5PHIB16 => return "L5PHIB16";
       when L5PHID31 => return "L5PHID31";
       when L4PHID29 => return "L4PHID29";
       when L4PHIA2 => return "L4PHIA2";
       when L5PHIB13 => return "L5PHIB13";
       when L1PHIG26 => return "L1PHIG26";
       when L3PHIB9 => return "L3PHIB9";
       when L2PHIB11 => return "L2PHIB11";
       when L3PHIC23 => return "L3PHIC23";
       when L3PHIA2 => return "L3PHIA2";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_AP_60) return string is
  begin
    case val is
       when L1PHIG => return "L1PHIG";
       when L1PHIA => return "L1PHIA";
       when L2PHID => return "L2PHID";
       when L3PHIB => return "L3PHIB";
       when L2PHIC => return "L2PHIC";
       when L3PHIC => return "L3PHIC";
       when L3PHIA => return "L3PHIA";
       when L1PHIH => return "L1PHIH";
       when L1PHIE => return "L1PHIE";
       when L1PHIF => return "L1PHIF";
       when L1PHID => return "L1PHID";
       when L3PHID => return "L3PHID";
       when L1PHIB => return "L1PHIB";
       when L2PHIB => return "L2PHIB";
       when L1PHIC => return "L1PHIC";
       when L2PHIA => return "L2PHIA";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_AP_58) return string is
  begin
    case val is
       when L4PHIA => return "L4PHIA";
       when L5PHIA => return "L5PHIA";
       when L5PHIB => return "L5PHIB";
       when L6PHIC => return "L6PHIC";
       when L6PHIB => return "L6PHIB";
       when L4PHIC => return "L4PHIC";
       when L4PHID => return "L4PHID";
       when L4PHIB => return "L4PHIB";
       when L6PHID => return "L6PHID";
       when L5PHIC => return "L5PHIC";
       when L6PHIA => return "L6PHIA";
       when L5PHID => return "L5PHID";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_CM_14) return string is
  begin
    case val is
       when L5PHIC17 => return "L5PHIC17";
       when L5PHIA5 => return "L5PHIA5";
       when L4PHID28 => return "L4PHID28";
       when L1PHID15 => return "L1PHID15";
       when L1PHIB6 => return "L1PHIB6";
       when L2PHID26 => return "L2PHID26";
       when L4PHID25 => return "L4PHID25";
       when L2PHIB15 => return "L2PHIB15";
       when L3PHIC20 => return "L3PHIC20";
       when L1PHIF22 => return "L1PHIF22";
       when L2PHIA4 => return "L2PHIA4";
       when L1PHIA1 => return "L1PHIA1";
       when L3PHIC23 => return "L3PHIC23";
       when L2PHID25 => return "L2PHID25";
       when L2PHID27 => return "L2PHID27";
       when L5PHIB13 => return "L5PHIB13";
       when L3PHIB9 => return "L3PHIB9";
       when L6PHIC18 => return "L6PHIC18";
       when L4PHIB11 => return "L4PHIB11";
       when L6PHIB15 => return "L6PHIB15";
       when L1PHIH29 => return "L1PHIH29";
       when L2PHID31 => return "L2PHID31";
       when L1PHID16 => return "L1PHID16";
       when L3PHID26 => return "L3PHID26";
       when L5PHIC24 => return "L5PHIC24";
       when L1PHIE17 => return "L1PHIE17";
       when L1PHIB7 => return "L1PHIB7";
       when L2PHID29 => return "L2PHID29";
       when L3PHIA4 => return "L3PHIA4";
       when L3PHIC22 => return "L3PHIC22";
       when L4PHIB14 => return "L4PHIB14";
       when L3PHID28 => return "L3PHID28";
       when L2PHIC23 => return "L2PHIC23";
       when L5PHID29 => return "L5PHID29";
       when L3PHIB12 => return "L3PHIB12";
       when L6PHIB13 => return "L6PHIB13";
       when L2PHIC21 => return "L2PHIC21";
       when L5PHIA6 => return "L5PHIA6";
       when L2PHIC19 => return "L2PHIC19";
       when L4PHIB12 => return "L4PHIB12";
       when L1PHIB5 => return "L1PHIB5";
       when L3PHIC24 => return "L3PHIC24";
       when L5PHIA7 => return "L5PHIA7";
       when L2PHIA3 => return "L2PHIA3";
       when L4PHID31 => return "L4PHID31";
       when L2PHIB12 => return "L2PHIB12";
       when L1PHIE18 => return "L1PHIE18";
       when L3PHIB11 => return "L3PHIB11";
       when L6PHIC20 => return "L6PHIC20";
       when L5PHIC20 => return "L5PHIC20";
       when L5PHID25 => return "L5PHID25";
       when L6PHIB11 => return "L6PHIB11";
       when L4PHIC17 => return "L4PHIC17";
       when L4PHIC21 => return "L4PHIC21";
       when L1PHIC11 => return "L1PHIC11";
       when L3PHIA2 => return "L3PHIA2";
       when L1PHID14 => return "L1PHID14";
       when L5PHIB14 => return "L5PHIB14";
       when L6PHID30 => return "L6PHID30";
       when L3PHIC18 => return "L3PHIC18";
       when L3PHID25 => return "L3PHID25";
       when L2PHID32 => return "L2PHID32";
       when L4PHIA7 => return "L4PHIA7";
       when L1PHIF21 => return "L1PHIF21";
       when L6PHIB10 => return "L6PHIB10";
       when L6PHIB9 => return "L6PHIB9";
       when L4PHIC22 => return "L4PHIC22";
       when L2PHIB10 => return "L2PHIB10";
       when L1PHID13 => return "L1PHID13";
       when L5PHIA2 => return "L5PHIA2";
       when L6PHIA7 => return "L6PHIA7";
       when L3PHIC21 => return "L3PHIC21";
       when L1PHIC12 => return "L1PHIC12";
       when L6PHID25 => return "L6PHID25";
       when L5PHIB16 => return "L5PHIB16";
       when L5PHID32 => return "L5PHID32";
       when L6PHID27 => return "L6PHID27";
       when L6PHIB12 => return "L6PHIB12";
       when L4PHIA6 => return "L4PHIA6";
       when L2PHIC22 => return "L2PHIC22";
       when L5PHIC19 => return "L5PHIC19";
       when L2PHIC18 => return "L2PHIC18";
       when L6PHIC24 => return "L6PHIC24";
       when L2PHIA2 => return "L2PHIA2";
       when L4PHIC19 => return "L4PHIC19";
       when L5PHIA3 => return "L5PHIA3";
       when L2PHIB13 => return "L2PHIB13";
       when L6PHIA8 => return "L6PHIA8";
       when L6PHID32 => return "L6PHID32";
       when L6PHIA2 => return "L6PHIA2";
       when L5PHIA4 => return "L5PHIA4";
       when L3PHIA8 => return "L3PHIA8";
       when L5PHIC21 => return "L5PHIC21";
       when L5PHIC18 => return "L5PHIC18";
       when L5PHIB9 => return "L5PHIB9";
       when L1PHIG26 => return "L1PHIG26";
       when L5PHIA1 => return "L5PHIA1";
       when L5PHID30 => return "L5PHID30";
       when L6PHIC23 => return "L6PHIC23";
       when L5PHIB10 => return "L5PHIB10";
       when L4PHIA5 => return "L4PHIA5";
       when L3PHIB14 => return "L3PHIB14";
       when L4PHID30 => return "L4PHID30";
       when L6PHIC19 => return "L6PHIC19";
       when L2PHIA1 => return "L2PHIA1";
       when L3PHIA6 => return "L3PHIA6";
       when L1PHIF24 => return "L1PHIF24";
       when L4PHIB10 => return "L4PHIB10";
       when L4PHIA8 => return "L4PHIA8";
       when L3PHID30 => return "L3PHID30";
       when L5PHIB12 => return "L5PHIB12";
       when L3PHID27 => return "L3PHID27";
       when L3PHIB10 => return "L3PHIB10";
       when L4PHIC20 => return "L4PHIC20";
       when L5PHID27 => return "L5PHID27";
       when L4PHID29 => return "L4PHID29";
       when L1PHIH30 => return "L1PHIH30";
       when L4PHIB16 => return "L4PHIB16";
       when L1PHIG28 => return "L1PHIG28";
       when L3PHIB13 => return "L3PHIB13";
       when L1PHIC9 => return "L1PHIC9";
       when L6PHIA1 => return "L6PHIA1";
       when L4PHID27 => return "L4PHID27";
       when L1PHIA4 => return "L1PHIA4";
       when L6PHID28 => return "L6PHID28";
       when L2PHIC24 => return "L2PHIC24";
       when L2PHIA7 => return "L2PHIA7";
       when L4PHIA4 => return "L4PHIA4";
       when L4PHIB15 => return "L4PHIB15";
       when L2PHIB14 => return "L2PHIB14";
       when L4PHIB13 => return "L4PHIB13";
       when L1PHIH31 => return "L1PHIH31";
       when L3PHIA7 => return "L3PHIA7";
       when L6PHID31 => return "L6PHID31";
       when L3PHIA1 => return "L3PHIA1";
       when L6PHID26 => return "L6PHID26";
       when L5PHIC22 => return "L5PHIC22";
       when L6PHIC21 => return "L6PHIC21";
       when L2PHIC17 => return "L2PHIC17";
       when L5PHID28 => return "L5PHID28";
       when L4PHIC24 => return "L4PHIC24";
       when L2PHIA6 => return "L2PHIA6";
       when L5PHIB11 => return "L5PHIB11";
       when L3PHIB16 => return "L3PHIB16";
       when L2PHIA8 => return "L2PHIA8";
       when L5PHID26 => return "L5PHID26";
       when L4PHID32 => return "L4PHID32";
       when L2PHIA5 => return "L2PHIA5";
       when L4PHID26 => return "L4PHID26";
       when L1PHIC10 => return "L1PHIC10";
       when L2PHID28 => return "L2PHID28";
       when L1PHIE20 => return "L1PHIE20";
       when L2PHID30 => return "L2PHID30";
       when L4PHIC18 => return "L4PHIC18";
       when L2PHIC20 => return "L2PHIC20";
       when L6PHIB14 => return "L6PHIB14";
       when L3PHID32 => return "L3PHID32";
       when L3PHIB15 => return "L3PHIB15";
       when L4PHIB9 => return "L4PHIB9";
       when L1PHIB8 => return "L1PHIB8";
       when L2PHIB9 => return "L2PHIB9";
       when L6PHIC22 => return "L6PHIC22";
       when L5PHIB15 => return "L5PHIB15";
       when L3PHIA3 => return "L3PHIA3";
       when L3PHID29 => return "L3PHID29";
       when L6PHIC17 => return "L6PHIC17";
       when L1PHIH32 => return "L1PHIH32";
       when L1PHIE19 => return "L1PHIE19";
       when L4PHIA3 => return "L4PHIA3";
       when L5PHID31 => return "L5PHID31";
       when L3PHIA5 => return "L3PHIA5";
       when L4PHIA1 => return "L4PHIA1";
       when L6PHID29 => return "L6PHID29";
       when L1PHIA2 => return "L1PHIA2";
       when L5PHIC23 => return "L5PHIC23";
       when L1PHIA3 => return "L1PHIA3";
       when L6PHIA4 => return "L6PHIA4";
       when L4PHIC23 => return "L4PHIC23";
       when L2PHIB16 => return "L2PHIB16";
       when L1PHIG25 => return "L1PHIG25";
       when L2PHIB11 => return "L2PHIB11";
       when L6PHIA3 => return "L6PHIA3";
       when L3PHIC19 => return "L3PHIC19";
       when L3PHID31 => return "L3PHID31";
       when L4PHIA2 => return "L4PHIA2";
       when L6PHIA5 => return "L6PHIA5";
       when L5PHIA8 => return "L5PHIA8";
       when L6PHIA6 => return "L6PHIA6";
       when L1PHIG27 => return "L1PHIG27";
       when L1PHIF23 => return "L1PHIF23";
       when L3PHIC17 => return "L3PHIC17";
       when L6PHIB16 => return "L6PHIB16";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_FM_52) return string is
  begin
    case val is
       when L5L6_L1PHIF => return "L5L6_L1PHIF";
       when L2L3_L1PHIG => return "L2L3_L1PHIG";
       when L2L3_L1PHID => return "L2L3_L1PHID";
       when L3L4_L5PHIB => return "L3L4_L5PHIB";
       when L3L4_L1PHIA => return "L3L4_L1PHIA";
       when L3L4_L1PHIC => return "L3L4_L1PHIC";
       when L1L2_L6PHIA => return "L1L2_L6PHIA";
       when L2L3_L5PHIB => return "L2L3_L5PHIB";
       when L2L3_L5PHIA => return "L2L3_L5PHIA";
       when L1L2_L3PHIA => return "L1L2_L3PHIA";
       when L3L4_L2PHID => return "L3L4_L2PHID";
       when L1L2_L5PHIC => return "L1L2_L5PHIC";
       when L2L3_L4PHIA => return "L2L3_L4PHIA";
       when L3L4_L1PHIH => return "L3L4_L1PHIH";
       when L5L6_L2PHIA => return "L5L6_L2PHIA";
       when L5L6_L3PHID => return "L5L6_L3PHID";
       when L3L4_L1PHIB => return "L3L4_L1PHIB";
       when L5L6_L4PHID => return "L5L6_L4PHID";
       when L1L2_L5PHIA => return "L1L2_L5PHIA";
       when L1L2_L4PHID => return "L1L2_L4PHID";
       when L2L3_L5PHID => return "L2L3_L5PHID";
       when L5L6_L2PHIB => return "L5L6_L2PHIB";
       when L1L2_L3PHID => return "L1L2_L3PHID";
       when L2L3_L4PHIB => return "L2L3_L4PHIB";
       when L1L2_L3PHIB => return "L1L2_L3PHIB";
       when L5L6_L3PHIA => return "L5L6_L3PHIA";
       when L2L3_L1PHIC => return "L2L3_L1PHIC";
       when L3L4_L1PHIF => return "L3L4_L1PHIF";
       when L3L4_L2PHIA => return "L3L4_L2PHIA";
       when L3L4_L6PHIB => return "L3L4_L6PHIB";
       when L2L3_L4PHID => return "L2L3_L4PHID";
       when L1L2_L4PHIB => return "L1L2_L4PHIB";
       when L3L4_L1PHID => return "L3L4_L1PHID";
       when L5L6_L1PHID => return "L5L6_L1PHID";
       when L3L4_L1PHIG => return "L3L4_L1PHIG";
       when L3L4_L1PHIE => return "L3L4_L1PHIE";
       when L2L3_L1PHIB => return "L2L3_L1PHIB";
       when L1L2_L3PHIC => return "L1L2_L3PHIC";
       when L2L3_L1PHIH => return "L2L3_L1PHIH";
       when L5L6_L4PHIC => return "L5L6_L4PHIC";
       when L3L4_L2PHIB => return "L3L4_L2PHIB";
       when L5L6_L1PHIG => return "L5L6_L1PHIG";
       when L1L2_L4PHIC => return "L1L2_L4PHIC";
       when L3L4_L2PHIC => return "L3L4_L2PHIC";
       when L2L3_L1PHIF => return "L2L3_L1PHIF";
       when L1L2_L4PHIA => return "L1L2_L4PHIA";
       when L3L4_L5PHIA => return "L3L4_L5PHIA";
       when L1L2_L5PHIB => return "L1L2_L5PHIB";
       when L5L6_L4PHIA => return "L5L6_L4PHIA";
       when L1L2_L6PHIC => return "L1L2_L6PHIC";
       when L3L4_L5PHID => return "L3L4_L5PHID";
       when L2L3_L1PHIA => return "L2L3_L1PHIA";
       when L1L2_L5PHID => return "L1L2_L5PHID";
       when L3L4_L6PHID => return "L3L4_L6PHID";
       when L5L6_L1PHIA => return "L5L6_L1PHIA";
       when L5L6_L3PHIC => return "L5L6_L3PHIC";
       when L1L2_L6PHIB => return "L1L2_L6PHIB";
       when L5L6_L1PHIH => return "L5L6_L1PHIH";
       when L5L6_L1PHIC => return "L5L6_L1PHIC";
       when L5L6_L1PHIB => return "L5L6_L1PHIB";
       when L3L4_L6PHIA => return "L3L4_L6PHIA";
       when L5L6_L1PHIE => return "L5L6_L1PHIE";
       when L3L4_L6PHIC => return "L3L4_L6PHIC";
       when L2L3_L1PHIE => return "L2L3_L1PHIE";
       when L5L6_L4PHIB => return "L5L6_L4PHIB";
       when L2L3_L4PHIC => return "L2L3_L4PHIC";
       when L3L4_L5PHIC => return "L3L4_L5PHIC";
       when L2L3_L5PHIC => return "L2L3_L5PHIC";
       when L5L6_L2PHID => return "L5L6_L2PHID";
       when L1L2_L6PHID => return "L1L2_L6PHID";
       when L5L6_L2PHIC => return "L5L6_L2PHIC";
       when L5L6_L3PHIB => return "L5L6_L3PHIB";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_TW_84) return string is
  begin
    case val is
       when L5L6 => return "L5L6";
       when L1L2 => return "L1L2";
       when L3L4 => return "L3L4";
       when L2L3 => return "L2L3";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

  function memory_enum_to_string(val: enum_BW_46) return string is
  begin
    case val is
       when L5L6_L1 => return "L5L6_L1";
       when L5L6_L2 => return "L5L6_L2";
       when L5L6_L3 => return "L5L6_L3";
       when L5L6_L4 => return "L5L6_L4";
       when L1L2_L3 => return "L1L2_L3";
       when L1L2_L4 => return "L1L2_L4";
       when L1L2_L5 => return "L1L2_L5";
       when L1L2_L6 => return "L1L2_L6";
       when L3L4_L1 => return "L3L4_L1";
       when L3L4_L2 => return "L3L4_L2";
       when L3L4_L5 => return "L3L4_L5";
       when L3L4_L6 => return "L3L4_L6";
       when L2L3_L1 => return "L2L3_L1";
       when L2L3_L4 => return "L2L3_L4";
       when L2L3_L5 => return "L2L3_L5";
    end case;
    return "No conversion found.";
  end memory_enum_to_string;

end package body memUtil_pkg;
