--! Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--! User packages
use work.tf_pkg.all;
use work.memUtil_pkg.all;

entity SectorProcessor is
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    TE_start  : in std_logic;
    TE_bx_in : in std_logic_vector(2 downto 0);
    TC_bx_out : out std_logic_vector(2 downto 0);
    TC_bx_out_vld : out std_logic;
    TC_done   : out std_logic;
    AS_36_mem_A_wea        : in t_arr_AS_36_1b;
    AS_36_mem_AV_writeaddr : in t_arr_AS_36_ADDR;
    AS_36_mem_AV_din       : in t_arr_AS_36_DATA;
    VMSTE_22_mem_A_wea        : in t_arr_VMSTE_22_1b;
    VMSTE_22_mem_AV_writeaddr : in t_arr_VMSTE_22_ADDR;
    VMSTE_22_mem_AV_din       : in t_arr_VMSTE_22_DATA;
    VMSTE_16_mem_A_wea        : in t_arr_VMSTE_16_1b;
    VMSTE_16_mem_AV_writeaddr : in t_arr_VMSTE_16_ADDR;
    VMSTE_16_mem_AV_din       : in t_arr_VMSTE_16_DATA;
    TPROJ_60_mem_A_enb          : in t_arr_TPROJ_60_1b;
    TPROJ_60_mem_AV_readaddr    : in t_arr_TPROJ_60_ADDR;
    TPROJ_60_mem_AV_dout        : out t_arr_TPROJ_60_DATA;
    TPROJ_60_mem_AAV_dout_nent  : out t_arr_TPROJ_60_NENT;
    TPROJ_58_mem_A_enb          : in t_arr_TPROJ_58_1b;
    TPROJ_58_mem_AV_readaddr    : in t_arr_TPROJ_58_ADDR;
    TPROJ_58_mem_AV_dout        : out t_arr_TPROJ_58_DATA;
    TPROJ_58_mem_AAV_dout_nent  : out t_arr_TPROJ_58_NENT;
    TPROJ_59_mem_A_enb          : in t_arr_TPROJ_59_1b;
    TPROJ_59_mem_AV_readaddr    : in t_arr_TPROJ_59_ADDR;
    TPROJ_59_mem_AV_dout        : out t_arr_TPROJ_59_DATA;
    TPROJ_59_mem_AAV_dout_nent  : out t_arr_TPROJ_59_NENT;
    TPAR_70_mem_A_enb          : in t_arr_TPAR_70_1b;
    TPAR_70_mem_AV_readaddr    : in t_arr_TPAR_70_ADDR;
    TPAR_70_mem_AV_dout        : out t_arr_TPAR_70_DATA;
    TPAR_70_mem_AAV_dout_nent  : out t_arr_TPAR_70_NENT
  );
end SectorProcessor;

architecture rtl of SectorProcessor is

  signal AS_36_mem_A_enb          : t_arr_AS_36_1b;
  signal AS_36_mem_AV_readaddr    : t_arr_AS_36_ADDR;
  signal AS_36_mem_AV_dout        : t_arr_AS_36_DATA;
  signal VMSTE_22_mem_A_enb          : t_arr_VMSTE_22_1b;
  signal VMSTE_22_mem_AV_readaddr    : t_arr_VMSTE_22_ADDR;
  signal VMSTE_22_mem_AV_dout        : t_arr_VMSTE_22_DATA;
  signal VMSTE_22_mem_AAV_dout_nent  : t_arr_VMSTE_22_NENT; -- (#page)
  signal VMSTE_16_mem_A_enb          : t_arr_VMSTE_16_1b;
  signal VMSTE_16_mem_AV_readaddr    : t_arr_VMSTE_16_ADDR;
  signal VMSTE_16_mem_AV_dout        : t_arr_VMSTE_16_DATA;
  signal VMSTE_16_mem_AAAV_dout_nent : t_arr_VMSTE_16_NENT; -- (#page)(#bin)
  signal SP_14_mem_A_wea          : t_arr_SP_14_1b;
  signal SP_14_mem_AV_writeaddr   : t_arr_SP_14_ADDR;
  signal SP_14_mem_AV_din         : t_arr_SP_14_DATA;
  signal SP_14_mem_A_enb          : t_arr_SP_14_1b;
  signal SP_14_mem_AV_readaddr    : t_arr_SP_14_ADDR;
  signal SP_14_mem_AV_dout        : t_arr_SP_14_DATA;
  signal SP_14_mem_AAV_dout_nent  : t_arr_SP_14_NENT; -- (#page)
  signal TPROJ_60_mem_A_wea          : t_arr_TPROJ_60_1b;
  signal TPROJ_60_mem_AV_writeaddr   : t_arr_TPROJ_60_ADDR;
  signal TPROJ_60_mem_AV_din         : t_arr_TPROJ_60_DATA;
  signal TPROJ_58_mem_A_wea          : t_arr_TPROJ_58_1b;
  signal TPROJ_58_mem_AV_writeaddr   : t_arr_TPROJ_58_ADDR;
  signal TPROJ_58_mem_AV_din         : t_arr_TPROJ_58_DATA;
  signal TPROJ_59_mem_A_wea          : t_arr_TPROJ_59_1b;
  signal TPROJ_59_mem_AV_writeaddr   : t_arr_TPROJ_59_ADDR;
  signal TPROJ_59_mem_AV_din         : t_arr_TPROJ_59_DATA;
  signal TPAR_70_mem_A_wea          : t_arr_TPAR_70_1b;
  signal TPAR_70_mem_AV_writeaddr   : t_arr_TPAR_70_ADDR;
  signal TPAR_70_mem_AV_din         : t_arr_TPAR_70_DATA;
  signal TE_done : std_logic := '0';
  signal TE_bx_out : std_logic_vector(2 downto 0);
  signal TE_bx_out_vld : std_logic;
  signal TC_start : std_logic := '0';
  signal TE_L1PHIC12_L2PHIB10_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB10_bendinnertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB10_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB10_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB10_bendoutertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB10_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB11_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB11_bendinnertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB11_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB11_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB11_bendoutertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB11_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB12_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB12_bendinnertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB12_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB12_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB12_bendoutertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB12_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB13_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB13_bendinnertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB13_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB13_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB13_bendoutertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB13_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB14_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB14_bendinnertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB14_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHIC12_L2PHIB14_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHIC12_L2PHIB14_bendoutertable_ce       : std_logic;
  signal TE_L1PHIC12_L2PHIB14_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB11_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB11_bendinnertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB11_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB11_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB11_bendoutertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB11_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB12_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB12_bendinnertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB12_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB12_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB12_bendoutertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB12_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB13_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB13_bendinnertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB13_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB13_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB13_bendoutertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB13_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB14_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB14_bendinnertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB14_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB14_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB14_bendoutertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB14_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB15_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB15_bendinnertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB15_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID13_L2PHIB15_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID13_L2PHIB15_bendoutertable_ce       : std_logic;
  signal TE_L1PHID13_L2PHIB15_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB12_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB12_bendinnertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB12_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB12_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB12_bendoutertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB12_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB13_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB13_bendinnertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB13_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB13_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB13_bendoutertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB13_bendoutertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB14_bendinnertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB14_bendinnertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB14_bendinnertable_dout : std_logic_vector(0 downto 0);
  signal TE_L1PHID14_L2PHIB14_bendoutertable_addr       : std_logic_vector(7 downto 0);
  signal TE_L1PHID14_L2PHIB14_bendoutertable_ce       : std_logic;
  signal TE_L1PHID14_L2PHIB14_bendoutertable_dout : std_logic_vector(0 downto 0);

begin

  AS_36_loop : for var in enum_AS_36 generate
  begin

    AS_36 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => AS_36_mem_A_wea(var),
        addra     => AS_36_mem_AV_writeaddr(var),
        dina      => AS_36_mem_AV_din(var),
        clkb      => clk,
        enb       => AS_36_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => AS_36_mem_AV_readaddr(var),
        doutb     => AS_36_mem_AV_dout(var),
        sync_nent => TC_start,
        nent_o    => open
      );

  end generate AS_36_loop;


  VMSTE_22_loop : for var in enum_VMSTE_22 generate
  begin

    VMSTE_22 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 22,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSTE_22_mem_A_wea(var),
        addra     => VMSTE_22_mem_AV_writeaddr(var),
        dina      => VMSTE_22_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSTE_22_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSTE_22_mem_AV_readaddr(var),
        doutb     => VMSTE_22_mem_AV_dout(var),
        sync_nent => TE_start,
        nent_o    => VMSTE_22_mem_AAV_dout_nent(var)
      );

  end generate VMSTE_22_loop;


  VMSTE_16_loop : for var in enum_VMSTE_16 generate
  begin

    VMSTE_16 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => VMSTE_16_mem_A_wea(var),
        addra     => VMSTE_16_mem_AV_writeaddr(var),
        dina      => VMSTE_16_mem_AV_din(var),
        clkb      => clk,
        enb       => VMSTE_16_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => VMSTE_16_mem_AV_readaddr(var),
        doutb     => VMSTE_16_mem_AV_dout(var),
        sync_nent => TE_start,
        nent_o    => VMSTE_16_mem_AAAV_dout_nent(var)
      );

  end generate VMSTE_16_loop;


  SP_14_loop : for var in enum_SP_14 generate
  begin

    SP_14 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 14,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => SP_14_mem_A_wea(var),
        addra     => SP_14_mem_AV_writeaddr(var),
        dina      => SP_14_mem_AV_din(var),
        clkb      => clk,
        enb       => SP_14_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => SP_14_mem_AV_readaddr(var),
        doutb     => SP_14_mem_AV_dout(var),
        sync_nent => TC_start,
        nent_o    => SP_14_mem_AAV_dout_nent(var)
      );

  end generate SP_14_loop;


  TPROJ_60_loop : for var in enum_TPROJ_60 generate
  begin

    TPROJ_60 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 60,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPROJ_60_mem_A_wea(var),
        addra     => TPROJ_60_mem_AV_writeaddr(var),
        dina      => TPROJ_60_mem_AV_din(var),
        clkb      => clk,
        enb       => TPROJ_60_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPROJ_60_mem_AV_readaddr(var),
        doutb     => TPROJ_60_mem_AV_dout(var),
        sync_nent => TC_done,
        nent_o    => TPROJ_60_mem_AAV_dout_nent(var)
      );

  end generate TPROJ_60_loop;


  TPROJ_58_loop : for var in enum_TPROJ_58 generate
  begin

    TPROJ_58 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 58,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPROJ_58_mem_A_wea(var),
        addra     => TPROJ_58_mem_AV_writeaddr(var),
        dina      => TPROJ_58_mem_AV_din(var),
        clkb      => clk,
        enb       => TPROJ_58_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPROJ_58_mem_AV_readaddr(var),
        doutb     => TPROJ_58_mem_AV_dout(var),
        sync_nent => TC_done,
        nent_o    => TPROJ_58_mem_AAV_dout_nent(var)
      );

  end generate TPROJ_58_loop;


  TPROJ_59_loop : for var in enum_TPROJ_59 generate
  begin

    TPROJ_59 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 59,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPROJ_59_mem_A_wea(var),
        addra     => TPROJ_59_mem_AV_writeaddr(var),
        dina      => TPROJ_59_mem_AV_din(var),
        clkb      => clk,
        enb       => TPROJ_59_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPROJ_59_mem_AV_readaddr(var),
        doutb     => TPROJ_59_mem_AV_dout(var),
        sync_nent => TC_done,
        nent_o    => TPROJ_59_mem_AAV_dout_nent(var)
      );

  end generate TPROJ_59_loop;


  TPAR_70_loop : for var in enum_TPAR_70 generate
  begin

    TPAR_70 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 70,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE"
      )
      port map (
        clka      => clk,
        wea       => TPAR_70_mem_A_wea(var),
        addra     => TPAR_70_mem_AV_writeaddr(var),
        dina      => TPAR_70_mem_AV_din(var),
        clkb      => clk,
        enb       => TPAR_70_mem_A_enb(var),
        rstb      => '0',
        regceb    => '1',
        addrb     => TPAR_70_mem_AV_readaddr(var),
        doutb     => TPAR_70_mem_AV_dout(var),
        sync_nent => TC_done,
        nent_o    => TPAR_70_mem_AAV_dout_nent(var)
      );

  end generate TPAR_70_loop;



  TE_L1PHIC12_L2PHIB10_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB10_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB10_bendinnertable_addr,
      ce        => TE_L1PHIC12_L2PHIB10_bendinnertable_ce,
      dout      => TE_L1PHIC12_L2PHIB10_bendinnertable_dout
  );


  TE_L1PHIC12_L2PHIB10_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB10_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB10_bendoutertable_addr,
      ce        => TE_L1PHIC12_L2PHIB10_bendoutertable_ce,
      dout      => TE_L1PHIC12_L2PHIB10_bendoutertable_dout
  );

  LATCH_TE: entity work.CreateStartSignal
    port map (
      clk   => clk,
      reset => reset,
      done  => TE_done,
      start => TC_start
  );

  TE_L1PHIC12_L2PHIB10 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TE_done,
      bx_V          => TE_bx_in,
      bx_o_V        => TE_bx_out,
      bx_o_V_ap_vld => TE_bx_out_vld,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHIC12n1),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHIC12n1),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHIC12n1),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n1)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n1)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB10n5),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB10n5),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB10n5),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB10n5)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHIC12_L2PHIB10_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHIC12_L2PHIB10_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHIC12_L2PHIB10_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHIC12_L2PHIB10_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHIC12_L2PHIB10_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHIC12_L2PHIB10_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHIC12_L2PHIB10),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHIC12_L2PHIB10),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHIC12_L2PHIB10)
  );


  TE_L1PHIC12_L2PHIB11_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB11_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB11_bendinnertable_addr,
      ce        => TE_L1PHIC12_L2PHIB11_bendinnertable_ce,
      dout      => TE_L1PHIC12_L2PHIB11_bendinnertable_dout
  );


  TE_L1PHIC12_L2PHIB11_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB11_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB11_bendoutertable_addr,
      ce        => TE_L1PHIC12_L2PHIB11_bendoutertable_ce,
      dout      => TE_L1PHIC12_L2PHIB11_bendoutertable_dout
  );

  TE_L1PHIC12_L2PHIB11 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHIC12n2),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHIC12n2),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHIC12n2),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n2)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n2)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB11n4),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB11n4),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB11n4),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n4)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHIC12_L2PHIB11_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHIC12_L2PHIB11_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHIC12_L2PHIB11_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHIC12_L2PHIB11_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHIC12_L2PHIB11_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHIC12_L2PHIB11_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHIC12_L2PHIB11),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHIC12_L2PHIB11),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHIC12_L2PHIB11)
  );


  TE_L1PHIC12_L2PHIB12_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB12_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB12_bendinnertable_addr,
      ce        => TE_L1PHIC12_L2PHIB12_bendinnertable_ce,
      dout      => TE_L1PHIC12_L2PHIB12_bendinnertable_dout
  );


  TE_L1PHIC12_L2PHIB12_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB12_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB12_bendoutertable_addr,
      ce        => TE_L1PHIC12_L2PHIB12_bendoutertable_ce,
      dout      => TE_L1PHIC12_L2PHIB12_bendoutertable_dout
  );

  TE_L1PHIC12_L2PHIB12 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHIC12n3),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHIC12n3),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHIC12n3),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n3)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n3)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB12n3),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB12n3),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB12n3),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n3)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHIC12_L2PHIB12_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHIC12_L2PHIB12_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHIC12_L2PHIB12_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHIC12_L2PHIB12_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHIC12_L2PHIB12_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHIC12_L2PHIB12_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHIC12_L2PHIB12),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHIC12_L2PHIB12),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHIC12_L2PHIB12)
  );


  TE_L1PHIC12_L2PHIB13_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB13_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB13_bendinnertable_addr,
      ce        => TE_L1PHIC12_L2PHIB13_bendinnertable_ce,
      dout      => TE_L1PHIC12_L2PHIB13_bendinnertable_dout
  );


  TE_L1PHIC12_L2PHIB13_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB13_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB13_bendoutertable_addr,
      ce        => TE_L1PHIC12_L2PHIB13_bendoutertable_ce,
      dout      => TE_L1PHIC12_L2PHIB13_bendoutertable_dout
  );

  TE_L1PHIC12_L2PHIB13 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHIC12n4),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHIC12n4),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHIC12n4),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n4)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n4)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB13n2),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB13n2),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB13n2),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n2)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHIC12_L2PHIB13_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHIC12_L2PHIB13_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHIC12_L2PHIB13_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHIC12_L2PHIB13_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHIC12_L2PHIB13_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHIC12_L2PHIB13_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHIC12_L2PHIB13),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHIC12_L2PHIB13),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHIC12_L2PHIB13)
  );


  TE_L1PHIC12_L2PHIB14_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB14_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB14_bendinnertable_addr,
      ce        => TE_L1PHIC12_L2PHIB14_bendinnertable_ce,
      dout      => TE_L1PHIC12_L2PHIB14_bendinnertable_dout
  );


  TE_L1PHIC12_L2PHIB14_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHIC12_L2PHIB14_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHIC12_L2PHIB14_bendoutertable_addr,
      ce        => TE_L1PHIC12_L2PHIB14_bendoutertable_ce,
      dout      => TE_L1PHIC12_L2PHIB14_bendoutertable_dout
  );

  TE_L1PHIC12_L2PHIB14 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHIC12n5),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHIC12n5),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHIC12n5),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n5)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHIC12n5)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB14n1),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB14n1),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB14n1),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n1)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHIC12_L2PHIB14_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHIC12_L2PHIB14_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHIC12_L2PHIB14_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHIC12_L2PHIB14_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHIC12_L2PHIB14_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHIC12_L2PHIB14_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHIC12_L2PHIB14),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHIC12_L2PHIB14),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHIC12_L2PHIB14)
  );


  TE_L1PHID13_L2PHIB11_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB11_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB11_bendinnertable_addr,
      ce        => TE_L1PHID13_L2PHIB11_bendinnertable_ce,
      dout      => TE_L1PHID13_L2PHIB11_bendinnertable_dout
  );


  TE_L1PHID13_L2PHIB11_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB11_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB11_bendoutertable_addr,
      ce        => TE_L1PHID13_L2PHIB11_bendoutertable_ce,
      dout      => TE_L1PHID13_L2PHIB11_bendoutertable_dout
  );

  TE_L1PHID13_L2PHIB11 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID13n1),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID13n1),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID13n1),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n1)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n1)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB11n5),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB11n5),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB11n5),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB11n5)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID13_L2PHIB11_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID13_L2PHIB11_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID13_L2PHIB11_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID13_L2PHIB11_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID13_L2PHIB11_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID13_L2PHIB11_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID13_L2PHIB11),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID13_L2PHIB11),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID13_L2PHIB11)
  );


  TE_L1PHID13_L2PHIB12_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB12_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB12_bendinnertable_addr,
      ce        => TE_L1PHID13_L2PHIB12_bendinnertable_ce,
      dout      => TE_L1PHID13_L2PHIB12_bendinnertable_dout
  );


  TE_L1PHID13_L2PHIB12_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB12_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB12_bendoutertable_addr,
      ce        => TE_L1PHID13_L2PHIB12_bendoutertable_ce,
      dout      => TE_L1PHID13_L2PHIB12_bendoutertable_dout
  );

  TE_L1PHID13_L2PHIB12 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID13n2),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID13n2),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID13n2),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n2)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n2)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB12n4),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB12n4),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB12n4),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n4)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID13_L2PHIB12_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID13_L2PHIB12_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID13_L2PHIB12_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID13_L2PHIB12_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID13_L2PHIB12_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID13_L2PHIB12_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID13_L2PHIB12),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID13_L2PHIB12),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID13_L2PHIB12)
  );


  TE_L1PHID13_L2PHIB13_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB13_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB13_bendinnertable_addr,
      ce        => TE_L1PHID13_L2PHIB13_bendinnertable_ce,
      dout      => TE_L1PHID13_L2PHIB13_bendinnertable_dout
  );


  TE_L1PHID13_L2PHIB13_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB13_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB13_bendoutertable_addr,
      ce        => TE_L1PHID13_L2PHIB13_bendoutertable_ce,
      dout      => TE_L1PHID13_L2PHIB13_bendoutertable_dout
  );

  TE_L1PHID13_L2PHIB13 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID13n3),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID13n3),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID13n3),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n3)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n3)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB13n3),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB13n3),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB13n3),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n3)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID13_L2PHIB13_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID13_L2PHIB13_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID13_L2PHIB13_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID13_L2PHIB13_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID13_L2PHIB13_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID13_L2PHIB13_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID13_L2PHIB13),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID13_L2PHIB13),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID13_L2PHIB13)
  );


  TE_L1PHID13_L2PHIB14_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB14_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB14_bendinnertable_addr,
      ce        => TE_L1PHID13_L2PHIB14_bendinnertable_ce,
      dout      => TE_L1PHID13_L2PHIB14_bendinnertable_dout
  );


  TE_L1PHID13_L2PHIB14_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB14_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB14_bendoutertable_addr,
      ce        => TE_L1PHID13_L2PHIB14_bendoutertable_ce,
      dout      => TE_L1PHID13_L2PHIB14_bendoutertable_dout
  );

  TE_L1PHID13_L2PHIB14 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID13n4),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID13n4),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID13n4),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n4)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n4)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB14n2),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB14n2),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB14n2),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n2)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID13_L2PHIB14_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID13_L2PHIB14_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID13_L2PHIB14_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID13_L2PHIB14_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID13_L2PHIB14_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID13_L2PHIB14_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID13_L2PHIB14),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID13_L2PHIB14),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID13_L2PHIB14)
  );


  TE_L1PHID13_L2PHIB15_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB15_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB15_bendinnertable_addr,
      ce        => TE_L1PHID13_L2PHIB15_bendinnertable_ce,
      dout      => TE_L1PHID13_L2PHIB15_bendinnertable_dout
  );


  TE_L1PHID13_L2PHIB15_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID13_L2PHIB15_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID13_L2PHIB15_bendoutertable_addr,
      ce        => TE_L1PHID13_L2PHIB15_bendoutertable_ce,
      dout      => TE_L1PHID13_L2PHIB15_bendoutertable_dout
  );

  TE_L1PHID13_L2PHIB15 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID13n5),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID13n5),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID13n5),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n5)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID13n5)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB15n1),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB15n1),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB15n1),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB15n1)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID13_L2PHIB15_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID13_L2PHIB15_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID13_L2PHIB15_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID13_L2PHIB15_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID13_L2PHIB15_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID13_L2PHIB15_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID13_L2PHIB15),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID13_L2PHIB15),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID13_L2PHIB15)
  );


  TE_L1PHID14_L2PHIB12_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB12_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB12_bendinnertable_addr,
      ce        => TE_L1PHID14_L2PHIB12_bendinnertable_ce,
      dout      => TE_L1PHID14_L2PHIB12_bendinnertable_dout
  );


  TE_L1PHID14_L2PHIB12_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB12_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB12_bendoutertable_addr,
      ce        => TE_L1PHID14_L2PHIB12_bendoutertable_ce,
      dout      => TE_L1PHID14_L2PHIB12_bendoutertable_dout
  );

  TE_L1PHID14_L2PHIB12 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID14n1),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID14n1),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID14n1),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n1)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n1)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB12n5),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB12n5),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB12n5),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB12n5)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID14_L2PHIB12_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID14_L2PHIB12_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID14_L2PHIB12_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID14_L2PHIB12_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID14_L2PHIB12_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID14_L2PHIB12_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID14_L2PHIB12),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID14_L2PHIB12),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID14_L2PHIB12)
  );


  TE_L1PHID14_L2PHIB13_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB13_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB13_bendinnertable_addr,
      ce        => TE_L1PHID14_L2PHIB13_bendinnertable_ce,
      dout      => TE_L1PHID14_L2PHIB13_bendinnertable_dout
  );


  TE_L1PHID14_L2PHIB13_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB13_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB13_bendoutertable_addr,
      ce        => TE_L1PHID14_L2PHIB13_bendoutertable_ce,
      dout      => TE_L1PHID14_L2PHIB13_bendoutertable_dout
  );

  TE_L1PHID14_L2PHIB13 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID14n2),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID14n2),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID14n2),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n2)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n2)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB13n4),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB13n4),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB13n4),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB13n4)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID14_L2PHIB13_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID14_L2PHIB13_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID14_L2PHIB13_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID14_L2PHIB13_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID14_L2PHIB13_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID14_L2PHIB13_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID14_L2PHIB13),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID14_L2PHIB13),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID14_L2PHIB13)
  );


  TE_L1PHID14_L2PHIB14_bendinnertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB14_stubptinnercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB14_bendinnertable_addr,
      ce        => TE_L1PHID14_L2PHIB14_bendinnertable_ce,
      dout      => TE_L1PHID14_L2PHIB14_bendinnertable_dout
  );


  TE_L1PHID14_L2PHIB14_bendoutertable : entity work.tf_lut
    generic map (
      lut_file  => "LUTs/TE_L1PHID14_L2PHIB14_stubptoutercut.tab",
      lut_width => 1,
      lut_depth => 256
    )
    port map (
      clk       => clk,
      addr      => TE_L1PHID14_L2PHIB14_bendoutertable_addr,
      ce        => TE_L1PHID14_L2PHIB14_bendoutertable_ce,
      dout      => TE_L1PHID14_L2PHIB14_bendoutertable_dout
  );

  TE_L1PHID14_L2PHIB14 : entity work.TE_L1L2
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TE_bx_in,
      instubinnerdata_dataarray_data_V_ce0       => VMSTE_22_mem_A_enb(L1PHID14n3),
      instubinnerdata_dataarray_data_V_address0  => VMSTE_22_mem_AV_readaddr(L1PHID14n3),
      instubinnerdata_dataarray_data_V_q0        => VMSTE_22_mem_AV_dout(L1PHID14n3),
      instubinnerdata_nentries_0_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n3)(0),
      instubinnerdata_nentries_1_V               => VMSTE_22_mem_AAV_dout_nent(L1PHID14n3)(1),
      instubouterdata_dataarray_data_V_ce0       => VMSTE_16_mem_A_enb(L2PHIB14n3),
      instubouterdata_dataarray_data_V_address0  => VMSTE_16_mem_AV_readaddr(L2PHIB14n3),
      instubouterdata_dataarray_data_V_q0        => VMSTE_16_mem_AV_dout(L2PHIB14n3),
      instubouterdata_nentries_0_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(0),
      instubouterdata_nentries_0_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(1),
      instubouterdata_nentries_0_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(2),
      instubouterdata_nentries_0_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(3),
      instubouterdata_nentries_0_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(4),
      instubouterdata_nentries_0_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(5),
      instubouterdata_nentries_0_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(6),
      instubouterdata_nentries_0_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(0)(7),
      instubouterdata_nentries_1_V_0     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(0),
      instubouterdata_nentries_1_V_1     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(1),
      instubouterdata_nentries_1_V_2     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(2),
      instubouterdata_nentries_1_V_3     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(3),
      instubouterdata_nentries_1_V_4     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(4),
      instubouterdata_nentries_1_V_5     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(5),
      instubouterdata_nentries_1_V_6     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(6),
      instubouterdata_nentries_1_V_7     => VMSTE_16_mem_AAAV_dout_nent(L2PHIB14n3)(1)(7),
      bendinnertable_V_address0                  => TE_L1PHID14_L2PHIB14_bendinnertable_addr,
      bendinnertable_V_ce0                       => TE_L1PHID14_L2PHIB14_bendinnertable_ce,
      bendinnertable_V_q0                        => TE_L1PHID14_L2PHIB14_bendinnertable_dout,
      bendoutertable_V_address0                  => TE_L1PHID14_L2PHIB14_bendoutertable_addr,
      bendoutertable_V_ce0                       => TE_L1PHID14_L2PHIB14_bendoutertable_ce,
      bendoutertable_V_q0                        => TE_L1PHID14_L2PHIB14_bendoutertable_dout,
      outstubpair_dataarray_data_V_ce0       => open,
      outstubpair_dataarray_data_V_we0       => SP_14_mem_A_wea(L1PHID14_L2PHIB14),
      outstubpair_dataarray_data_V_address0  => SP_14_mem_AV_writeaddr(L1PHID14_L2PHIB14),
      outstubpair_dataarray_data_V_d0        => SP_14_mem_AV_din(L1PHID14_L2PHIB14)
  );

  TC_L1L2E : entity work.TC_L1L2E
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TC_done,
      bx_V          => TE_bx_out,
      bx_o_V        => TC_bx_out,
      bx_o_V_ap_vld => TC_bx_out_vld,
      innerStubs_0_dataarray_data_V_ce0       => AS_36_mem_A_enb(L1PHICn4),
      innerStubs_0_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L1PHICn4),
      innerStubs_0_dataarray_data_V_q0        => AS_36_mem_AV_dout(L1PHICn4),
      innerStubs_1_dataarray_data_V_ce0       => AS_36_mem_A_enb(L1PHIDn2),
      innerStubs_1_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L1PHIDn2),
      innerStubs_1_dataarray_data_V_q0        => AS_36_mem_AV_dout(L1PHIDn2),
      outerStubs_0_dataarray_data_V_ce0       => AS_36_mem_A_enb(L2PHIBn4),
      outerStubs_0_dataarray_data_V_address0  => AS_36_mem_AV_readaddr(L2PHIBn4),
      outerStubs_0_dataarray_data_V_q0        => AS_36_mem_AV_dout(L2PHIBn4),
      stubPairs_0_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHIC12_L2PHIB10),
      stubPairs_0_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHIC12_L2PHIB10),
      stubPairs_0_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHIC12_L2PHIB10),
      stubPairs_0_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB10)(0),
      stubPairs_0_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB10)(1),
      stubPairs_1_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHIC12_L2PHIB11),
      stubPairs_1_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHIC12_L2PHIB11),
      stubPairs_1_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHIC12_L2PHIB11),
      stubPairs_1_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB11)(0),
      stubPairs_1_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB11)(1),
      stubPairs_2_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHIC12_L2PHIB12),
      stubPairs_2_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHIC12_L2PHIB12),
      stubPairs_2_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHIC12_L2PHIB12),
      stubPairs_2_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB12)(0),
      stubPairs_2_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB12)(1),
      stubPairs_3_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHIC12_L2PHIB13),
      stubPairs_3_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHIC12_L2PHIB13),
      stubPairs_3_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHIC12_L2PHIB13),
      stubPairs_3_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB13)(0),
      stubPairs_3_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB13)(1),
      stubPairs_4_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHIC12_L2PHIB14),
      stubPairs_4_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHIC12_L2PHIB14),
      stubPairs_4_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHIC12_L2PHIB14),
      stubPairs_4_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB14)(0),
      stubPairs_4_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHIC12_L2PHIB14)(1),
      stubPairs_5_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID13_L2PHIB11),
      stubPairs_5_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID13_L2PHIB11),
      stubPairs_5_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID13_L2PHIB11),
      stubPairs_5_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB11)(0),
      stubPairs_5_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB11)(1),
      stubPairs_6_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID13_L2PHIB12),
      stubPairs_6_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID13_L2PHIB12),
      stubPairs_6_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID13_L2PHIB12),
      stubPairs_6_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB12)(0),
      stubPairs_6_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB12)(1),
      stubPairs_7_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID13_L2PHIB13),
      stubPairs_7_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID13_L2PHIB13),
      stubPairs_7_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID13_L2PHIB13),
      stubPairs_7_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB13)(0),
      stubPairs_7_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB13)(1),
      stubPairs_8_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID13_L2PHIB14),
      stubPairs_8_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID13_L2PHIB14),
      stubPairs_8_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID13_L2PHIB14),
      stubPairs_8_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB14)(0),
      stubPairs_8_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB14)(1),
      stubPairs_9_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID13_L2PHIB15),
      stubPairs_9_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID13_L2PHIB15),
      stubPairs_9_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID13_L2PHIB15),
      stubPairs_9_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB15)(0),
      stubPairs_9_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID13_L2PHIB15)(1),
      stubPairs_10_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID14_L2PHIB12),
      stubPairs_10_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID14_L2PHIB12),
      stubPairs_10_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID14_L2PHIB12),
      stubPairs_10_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB12)(0),
      stubPairs_10_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB12)(1),
      stubPairs_11_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID14_L2PHIB13),
      stubPairs_11_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID14_L2PHIB13),
      stubPairs_11_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID14_L2PHIB13),
      stubPairs_11_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB13)(0),
      stubPairs_11_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB13)(1),
      stubPairs_12_dataarray_data_V_ce0       => SP_14_mem_A_enb(L1PHID14_L2PHIB14),
      stubPairs_12_dataarray_data_V_address0  => SP_14_mem_AV_readaddr(L1PHID14_L2PHIB14),
      stubPairs_12_dataarray_data_V_q0        => SP_14_mem_AV_dout(L1PHID14_L2PHIB14),
      stubPairs_12_nentries_0_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB14)(0),
      stubPairs_12_nentries_1_V               => SP_14_mem_AAV_dout_nent(L1PHID14_L2PHIB14)(1),
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_70_mem_A_wea(L1L2E),
      trackletParameters_dataarray_data_V_address0  => TPAR_70_mem_AV_writeaddr(L1L2E),
      trackletParameters_dataarray_data_V_d0        => TPAR_70_mem_AV_din(L1L2E),
      projout_barrel_ps_13_dataarray_data_V_ce0       => open,
      projout_barrel_ps_13_dataarray_data_V_we0       => TPROJ_60_mem_A_wea(L1L2E_L3PHIB),
      projout_barrel_ps_13_dataarray_data_V_address0  => TPROJ_60_mem_AV_writeaddr(L1L2E_L3PHIB),
      projout_barrel_ps_13_dataarray_data_V_d0        => TPROJ_60_mem_AV_din(L1L2E_L3PHIB),
      projout_barrel_2s_0_dataarray_data_V_ce0       => open,
      projout_barrel_2s_0_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L4PHIA),
      projout_barrel_2s_0_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L4PHIA),
      projout_barrel_2s_0_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L4PHIA),
      projout_barrel_2s_1_dataarray_data_V_ce0       => open,
      projout_barrel_2s_1_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L4PHIB),
      projout_barrel_2s_1_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L4PHIB),
      projout_barrel_2s_1_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L4PHIB),
      projout_barrel_2s_2_dataarray_data_V_ce0       => open,
      projout_barrel_2s_2_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L4PHIC),
      projout_barrel_2s_2_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L4PHIC),
      projout_barrel_2s_2_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L4PHIC),
      projout_barrel_2s_4_dataarray_data_V_ce0       => open,
      projout_barrel_2s_4_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L5PHIA),
      projout_barrel_2s_4_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L5PHIA),
      projout_barrel_2s_4_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L5PHIA),
      projout_barrel_2s_5_dataarray_data_V_ce0       => open,
      projout_barrel_2s_5_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L5PHIB),
      projout_barrel_2s_5_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L5PHIB),
      projout_barrel_2s_5_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L5PHIB),
      projout_barrel_2s_6_dataarray_data_V_ce0       => open,
      projout_barrel_2s_6_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L5PHIC),
      projout_barrel_2s_6_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L5PHIC),
      projout_barrel_2s_6_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L5PHIC),
      projout_barrel_2s_8_dataarray_data_V_ce0       => open,
      projout_barrel_2s_8_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L6PHIA),
      projout_barrel_2s_8_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L6PHIA),
      projout_barrel_2s_8_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L6PHIA),
      projout_barrel_2s_9_dataarray_data_V_ce0       => open,
      projout_barrel_2s_9_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L6PHIB),
      projout_barrel_2s_9_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L6PHIB),
      projout_barrel_2s_9_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L6PHIB),
      projout_barrel_2s_10_dataarray_data_V_ce0       => open,
      projout_barrel_2s_10_dataarray_data_V_we0       => TPROJ_58_mem_A_wea(L1L2E_L6PHIC),
      projout_barrel_2s_10_dataarray_data_V_address0  => TPROJ_58_mem_AV_writeaddr(L1L2E_L6PHIC),
      projout_barrel_2s_10_dataarray_data_V_d0        => TPROJ_58_mem_AV_din(L1L2E_L6PHIC),
      projout_disk_0_dataarray_data_V_ce0       => open,
      projout_disk_0_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D1PHIA),
      projout_disk_0_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D1PHIA),
      projout_disk_0_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D1PHIA),
      projout_disk_1_dataarray_data_V_ce0       => open,
      projout_disk_1_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D1PHIB),
      projout_disk_1_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D1PHIB),
      projout_disk_1_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D1PHIB),
      projout_disk_2_dataarray_data_V_ce0       => open,
      projout_disk_2_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D1PHIC),
      projout_disk_2_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D1PHIC),
      projout_disk_2_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D1PHIC),
      projout_disk_4_dataarray_data_V_ce0       => open,
      projout_disk_4_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D2PHIA),
      projout_disk_4_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D2PHIA),
      projout_disk_4_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D2PHIA),
      projout_disk_5_dataarray_data_V_ce0       => open,
      projout_disk_5_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D2PHIB),
      projout_disk_5_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D2PHIB),
      projout_disk_5_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D2PHIB),
      projout_disk_6_dataarray_data_V_ce0       => open,
      projout_disk_6_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D2PHIC),
      projout_disk_6_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D2PHIC),
      projout_disk_6_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D2PHIC),
      projout_disk_8_dataarray_data_V_ce0       => open,
      projout_disk_8_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D3PHIA),
      projout_disk_8_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D3PHIA),
      projout_disk_8_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D3PHIA),
      projout_disk_9_dataarray_data_V_ce0       => open,
      projout_disk_9_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D3PHIB),
      projout_disk_9_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D3PHIB),
      projout_disk_9_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D3PHIB),
      projout_disk_10_dataarray_data_V_ce0       => open,
      projout_disk_10_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D3PHIC),
      projout_disk_10_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D3PHIC),
      projout_disk_10_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D3PHIC),
      projout_disk_12_dataarray_data_V_ce0       => open,
      projout_disk_12_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D4PHIA),
      projout_disk_12_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D4PHIA),
      projout_disk_12_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D4PHIA),
      projout_disk_13_dataarray_data_V_ce0       => open,
      projout_disk_13_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D4PHIB),
      projout_disk_13_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D4PHIB),
      projout_disk_13_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D4PHIB),
      projout_disk_14_dataarray_data_V_ce0       => open,
      projout_disk_14_dataarray_data_V_we0       => TPROJ_59_mem_A_wea(L1L2E_D4PHIC),
      projout_disk_14_dataarray_data_V_address0  => TPROJ_59_mem_AV_writeaddr(L1L2E_D4PHIC),
      projout_disk_14_dataarray_data_V_d0        => TPROJ_59_mem_AV_din(L1L2E_D4PHIC)
  );



end rtl;
